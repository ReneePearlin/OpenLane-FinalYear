module picorv32_wrapper (clk,
    mem_instr,
    mem_ready,
    mem_valid,
    resetn,
    trap,
    mem_addr,
    mem_rdata,
    mem_wdata,
    mem_wstrb);
 input clk;
 output mem_instr;
 input mem_ready;
 output mem_valid;
 input resetn;
 output trap;
 output [31:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire \core.alu_out[0] ;
 wire \core.alu_out[10] ;
 wire \core.alu_out[11] ;
 wire \core.alu_out[12] ;
 wire \core.alu_out[13] ;
 wire \core.alu_out[14] ;
 wire \core.alu_out[15] ;
 wire \core.alu_out[16] ;
 wire \core.alu_out[17] ;
 wire \core.alu_out[18] ;
 wire \core.alu_out[19] ;
 wire \core.alu_out[1] ;
 wire \core.alu_out[20] ;
 wire \core.alu_out[21] ;
 wire \core.alu_out[22] ;
 wire \core.alu_out[23] ;
 wire \core.alu_out[24] ;
 wire \core.alu_out[25] ;
 wire \core.alu_out[26] ;
 wire \core.alu_out[27] ;
 wire \core.alu_out[28] ;
 wire \core.alu_out[29] ;
 wire \core.alu_out[2] ;
 wire \core.alu_out[30] ;
 wire \core.alu_out[31] ;
 wire \core.alu_out[3] ;
 wire \core.alu_out[4] ;
 wire \core.alu_out[5] ;
 wire \core.alu_out[6] ;
 wire \core.alu_out[7] ;
 wire \core.alu_out[8] ;
 wire \core.alu_out[9] ;
 wire \core.alu_out_q[0] ;
 wire \core.alu_out_q[10] ;
 wire \core.alu_out_q[11] ;
 wire \core.alu_out_q[12] ;
 wire \core.alu_out_q[13] ;
 wire \core.alu_out_q[14] ;
 wire \core.alu_out_q[15] ;
 wire \core.alu_out_q[16] ;
 wire \core.alu_out_q[17] ;
 wire \core.alu_out_q[18] ;
 wire \core.alu_out_q[19] ;
 wire \core.alu_out_q[1] ;
 wire \core.alu_out_q[20] ;
 wire \core.alu_out_q[21] ;
 wire \core.alu_out_q[22] ;
 wire \core.alu_out_q[23] ;
 wire \core.alu_out_q[24] ;
 wire \core.alu_out_q[25] ;
 wire \core.alu_out_q[26] ;
 wire \core.alu_out_q[27] ;
 wire \core.alu_out_q[28] ;
 wire \core.alu_out_q[29] ;
 wire \core.alu_out_q[2] ;
 wire \core.alu_out_q[30] ;
 wire \core.alu_out_q[31] ;
 wire \core.alu_out_q[3] ;
 wire \core.alu_out_q[4] ;
 wire \core.alu_out_q[5] ;
 wire \core.alu_out_q[6] ;
 wire \core.alu_out_q[7] ;
 wire \core.alu_out_q[8] ;
 wire \core.alu_out_q[9] ;
 wire \core.count_cycle[0] ;
 wire \core.count_cycle[10] ;
 wire \core.count_cycle[11] ;
 wire \core.count_cycle[12] ;
 wire \core.count_cycle[13] ;
 wire \core.count_cycle[14] ;
 wire \core.count_cycle[15] ;
 wire \core.count_cycle[16] ;
 wire \core.count_cycle[17] ;
 wire \core.count_cycle[18] ;
 wire \core.count_cycle[19] ;
 wire \core.count_cycle[1] ;
 wire \core.count_cycle[20] ;
 wire \core.count_cycle[21] ;
 wire \core.count_cycle[22] ;
 wire \core.count_cycle[23] ;
 wire \core.count_cycle[24] ;
 wire \core.count_cycle[25] ;
 wire \core.count_cycle[26] ;
 wire \core.count_cycle[27] ;
 wire \core.count_cycle[28] ;
 wire \core.count_cycle[29] ;
 wire \core.count_cycle[2] ;
 wire \core.count_cycle[30] ;
 wire \core.count_cycle[31] ;
 wire \core.count_cycle[32] ;
 wire \core.count_cycle[33] ;
 wire \core.count_cycle[34] ;
 wire \core.count_cycle[35] ;
 wire \core.count_cycle[36] ;
 wire \core.count_cycle[37] ;
 wire \core.count_cycle[38] ;
 wire \core.count_cycle[39] ;
 wire \core.count_cycle[3] ;
 wire \core.count_cycle[40] ;
 wire \core.count_cycle[41] ;
 wire \core.count_cycle[42] ;
 wire \core.count_cycle[43] ;
 wire \core.count_cycle[44] ;
 wire \core.count_cycle[45] ;
 wire \core.count_cycle[46] ;
 wire \core.count_cycle[47] ;
 wire \core.count_cycle[48] ;
 wire \core.count_cycle[49] ;
 wire \core.count_cycle[4] ;
 wire \core.count_cycle[50] ;
 wire \core.count_cycle[51] ;
 wire \core.count_cycle[52] ;
 wire \core.count_cycle[53] ;
 wire \core.count_cycle[54] ;
 wire \core.count_cycle[55] ;
 wire \core.count_cycle[56] ;
 wire \core.count_cycle[57] ;
 wire \core.count_cycle[58] ;
 wire \core.count_cycle[59] ;
 wire \core.count_cycle[5] ;
 wire \core.count_cycle[60] ;
 wire \core.count_cycle[61] ;
 wire \core.count_cycle[62] ;
 wire \core.count_cycle[63] ;
 wire \core.count_cycle[6] ;
 wire \core.count_cycle[7] ;
 wire \core.count_cycle[8] ;
 wire \core.count_cycle[9] ;
 wire \core.count_instr[0] ;
 wire \core.count_instr[10] ;
 wire \core.count_instr[11] ;
 wire \core.count_instr[12] ;
 wire \core.count_instr[13] ;
 wire \core.count_instr[14] ;
 wire \core.count_instr[15] ;
 wire \core.count_instr[16] ;
 wire \core.count_instr[17] ;
 wire \core.count_instr[18] ;
 wire \core.count_instr[19] ;
 wire \core.count_instr[1] ;
 wire \core.count_instr[20] ;
 wire \core.count_instr[21] ;
 wire \core.count_instr[22] ;
 wire \core.count_instr[23] ;
 wire \core.count_instr[24] ;
 wire \core.count_instr[25] ;
 wire \core.count_instr[26] ;
 wire \core.count_instr[27] ;
 wire \core.count_instr[28] ;
 wire \core.count_instr[29] ;
 wire \core.count_instr[2] ;
 wire \core.count_instr[30] ;
 wire \core.count_instr[31] ;
 wire \core.count_instr[32] ;
 wire \core.count_instr[33] ;
 wire \core.count_instr[34] ;
 wire \core.count_instr[35] ;
 wire \core.count_instr[36] ;
 wire \core.count_instr[37] ;
 wire \core.count_instr[38] ;
 wire \core.count_instr[39] ;
 wire \core.count_instr[3] ;
 wire \core.count_instr[40] ;
 wire \core.count_instr[41] ;
 wire \core.count_instr[42] ;
 wire \core.count_instr[43] ;
 wire \core.count_instr[44] ;
 wire \core.count_instr[45] ;
 wire \core.count_instr[46] ;
 wire \core.count_instr[47] ;
 wire \core.count_instr[48] ;
 wire \core.count_instr[49] ;
 wire \core.count_instr[4] ;
 wire \core.count_instr[50] ;
 wire \core.count_instr[51] ;
 wire \core.count_instr[52] ;
 wire \core.count_instr[53] ;
 wire \core.count_instr[54] ;
 wire \core.count_instr[55] ;
 wire \core.count_instr[56] ;
 wire \core.count_instr[57] ;
 wire \core.count_instr[58] ;
 wire \core.count_instr[59] ;
 wire \core.count_instr[5] ;
 wire \core.count_instr[60] ;
 wire \core.count_instr[61] ;
 wire \core.count_instr[62] ;
 wire \core.count_instr[63] ;
 wire \core.count_instr[6] ;
 wire \core.count_instr[7] ;
 wire \core.count_instr[8] ;
 wire \core.count_instr[9] ;
 wire \core.cpu_state[0] ;
 wire \core.cpu_state[1] ;
 wire \core.cpu_state[2] ;
 wire \core.cpu_state[3] ;
 wire \core.cpu_state[4] ;
 wire \core.cpu_state[5] ;
 wire \core.cpu_state[6] ;
 wire \core.cpuregs[0][0] ;
 wire \core.cpuregs[0][10] ;
 wire \core.cpuregs[0][11] ;
 wire \core.cpuregs[0][12] ;
 wire \core.cpuregs[0][13] ;
 wire \core.cpuregs[0][14] ;
 wire \core.cpuregs[0][15] ;
 wire \core.cpuregs[0][16] ;
 wire \core.cpuregs[0][17] ;
 wire \core.cpuregs[0][18] ;
 wire \core.cpuregs[0][19] ;
 wire \core.cpuregs[0][1] ;
 wire \core.cpuregs[0][20] ;
 wire \core.cpuregs[0][21] ;
 wire \core.cpuregs[0][22] ;
 wire \core.cpuregs[0][23] ;
 wire \core.cpuregs[0][24] ;
 wire \core.cpuregs[0][25] ;
 wire \core.cpuregs[0][26] ;
 wire \core.cpuregs[0][27] ;
 wire \core.cpuregs[0][28] ;
 wire \core.cpuregs[0][29] ;
 wire \core.cpuregs[0][2] ;
 wire \core.cpuregs[0][30] ;
 wire \core.cpuregs[0][31] ;
 wire \core.cpuregs[0][3] ;
 wire \core.cpuregs[0][4] ;
 wire \core.cpuregs[0][5] ;
 wire \core.cpuregs[0][6] ;
 wire \core.cpuregs[0][7] ;
 wire \core.cpuregs[0][8] ;
 wire \core.cpuregs[0][9] ;
 wire \core.cpuregs[10][0] ;
 wire \core.cpuregs[10][10] ;
 wire \core.cpuregs[10][11] ;
 wire \core.cpuregs[10][12] ;
 wire \core.cpuregs[10][13] ;
 wire \core.cpuregs[10][14] ;
 wire \core.cpuregs[10][15] ;
 wire \core.cpuregs[10][16] ;
 wire \core.cpuregs[10][17] ;
 wire \core.cpuregs[10][18] ;
 wire \core.cpuregs[10][19] ;
 wire \core.cpuregs[10][1] ;
 wire \core.cpuregs[10][20] ;
 wire \core.cpuregs[10][21] ;
 wire \core.cpuregs[10][22] ;
 wire \core.cpuregs[10][23] ;
 wire \core.cpuregs[10][24] ;
 wire \core.cpuregs[10][25] ;
 wire \core.cpuregs[10][26] ;
 wire \core.cpuregs[10][27] ;
 wire \core.cpuregs[10][28] ;
 wire \core.cpuregs[10][29] ;
 wire \core.cpuregs[10][2] ;
 wire \core.cpuregs[10][30] ;
 wire \core.cpuregs[10][31] ;
 wire \core.cpuregs[10][3] ;
 wire \core.cpuregs[10][4] ;
 wire \core.cpuregs[10][5] ;
 wire \core.cpuregs[10][6] ;
 wire \core.cpuregs[10][7] ;
 wire \core.cpuregs[10][8] ;
 wire \core.cpuregs[10][9] ;
 wire \core.cpuregs[11][0] ;
 wire \core.cpuregs[11][10] ;
 wire \core.cpuregs[11][11] ;
 wire \core.cpuregs[11][12] ;
 wire \core.cpuregs[11][13] ;
 wire \core.cpuregs[11][14] ;
 wire \core.cpuregs[11][15] ;
 wire \core.cpuregs[11][16] ;
 wire \core.cpuregs[11][17] ;
 wire \core.cpuregs[11][18] ;
 wire \core.cpuregs[11][19] ;
 wire \core.cpuregs[11][1] ;
 wire \core.cpuregs[11][20] ;
 wire \core.cpuregs[11][21] ;
 wire \core.cpuregs[11][22] ;
 wire \core.cpuregs[11][23] ;
 wire \core.cpuregs[11][24] ;
 wire \core.cpuregs[11][25] ;
 wire \core.cpuregs[11][26] ;
 wire \core.cpuregs[11][27] ;
 wire \core.cpuregs[11][28] ;
 wire \core.cpuregs[11][29] ;
 wire \core.cpuregs[11][2] ;
 wire \core.cpuregs[11][30] ;
 wire \core.cpuregs[11][31] ;
 wire \core.cpuregs[11][3] ;
 wire \core.cpuregs[11][4] ;
 wire \core.cpuregs[11][5] ;
 wire \core.cpuregs[11][6] ;
 wire \core.cpuregs[11][7] ;
 wire \core.cpuregs[11][8] ;
 wire \core.cpuregs[11][9] ;
 wire \core.cpuregs[12][0] ;
 wire \core.cpuregs[12][10] ;
 wire \core.cpuregs[12][11] ;
 wire \core.cpuregs[12][12] ;
 wire \core.cpuregs[12][13] ;
 wire \core.cpuregs[12][14] ;
 wire \core.cpuregs[12][15] ;
 wire \core.cpuregs[12][16] ;
 wire \core.cpuregs[12][17] ;
 wire \core.cpuregs[12][18] ;
 wire \core.cpuregs[12][19] ;
 wire \core.cpuregs[12][1] ;
 wire \core.cpuregs[12][20] ;
 wire \core.cpuregs[12][21] ;
 wire \core.cpuregs[12][22] ;
 wire \core.cpuregs[12][23] ;
 wire \core.cpuregs[12][24] ;
 wire \core.cpuregs[12][25] ;
 wire \core.cpuregs[12][26] ;
 wire \core.cpuregs[12][27] ;
 wire \core.cpuregs[12][28] ;
 wire \core.cpuregs[12][29] ;
 wire \core.cpuregs[12][2] ;
 wire \core.cpuregs[12][30] ;
 wire \core.cpuregs[12][31] ;
 wire \core.cpuregs[12][3] ;
 wire \core.cpuregs[12][4] ;
 wire \core.cpuregs[12][5] ;
 wire \core.cpuregs[12][6] ;
 wire \core.cpuregs[12][7] ;
 wire \core.cpuregs[12][8] ;
 wire \core.cpuregs[12][9] ;
 wire \core.cpuregs[13][0] ;
 wire \core.cpuregs[13][10] ;
 wire \core.cpuregs[13][11] ;
 wire \core.cpuregs[13][12] ;
 wire \core.cpuregs[13][13] ;
 wire \core.cpuregs[13][14] ;
 wire \core.cpuregs[13][15] ;
 wire \core.cpuregs[13][16] ;
 wire \core.cpuregs[13][17] ;
 wire \core.cpuregs[13][18] ;
 wire \core.cpuregs[13][19] ;
 wire \core.cpuregs[13][1] ;
 wire \core.cpuregs[13][20] ;
 wire \core.cpuregs[13][21] ;
 wire \core.cpuregs[13][22] ;
 wire \core.cpuregs[13][23] ;
 wire \core.cpuregs[13][24] ;
 wire \core.cpuregs[13][25] ;
 wire \core.cpuregs[13][26] ;
 wire \core.cpuregs[13][27] ;
 wire \core.cpuregs[13][28] ;
 wire \core.cpuregs[13][29] ;
 wire \core.cpuregs[13][2] ;
 wire \core.cpuregs[13][30] ;
 wire \core.cpuregs[13][31] ;
 wire \core.cpuregs[13][3] ;
 wire \core.cpuregs[13][4] ;
 wire \core.cpuregs[13][5] ;
 wire \core.cpuregs[13][6] ;
 wire \core.cpuregs[13][7] ;
 wire \core.cpuregs[13][8] ;
 wire \core.cpuregs[13][9] ;
 wire \core.cpuregs[14][0] ;
 wire \core.cpuregs[14][10] ;
 wire \core.cpuregs[14][11] ;
 wire \core.cpuregs[14][12] ;
 wire \core.cpuregs[14][13] ;
 wire \core.cpuregs[14][14] ;
 wire \core.cpuregs[14][15] ;
 wire \core.cpuregs[14][16] ;
 wire \core.cpuregs[14][17] ;
 wire \core.cpuregs[14][18] ;
 wire \core.cpuregs[14][19] ;
 wire \core.cpuregs[14][1] ;
 wire \core.cpuregs[14][20] ;
 wire \core.cpuregs[14][21] ;
 wire \core.cpuregs[14][22] ;
 wire \core.cpuregs[14][23] ;
 wire \core.cpuregs[14][24] ;
 wire \core.cpuregs[14][25] ;
 wire \core.cpuregs[14][26] ;
 wire \core.cpuregs[14][27] ;
 wire \core.cpuregs[14][28] ;
 wire \core.cpuregs[14][29] ;
 wire \core.cpuregs[14][2] ;
 wire \core.cpuregs[14][30] ;
 wire \core.cpuregs[14][31] ;
 wire \core.cpuregs[14][3] ;
 wire \core.cpuregs[14][4] ;
 wire \core.cpuregs[14][5] ;
 wire \core.cpuregs[14][6] ;
 wire \core.cpuregs[14][7] ;
 wire \core.cpuregs[14][8] ;
 wire \core.cpuregs[14][9] ;
 wire \core.cpuregs[15][0] ;
 wire \core.cpuregs[15][10] ;
 wire \core.cpuregs[15][11] ;
 wire \core.cpuregs[15][12] ;
 wire \core.cpuregs[15][13] ;
 wire \core.cpuregs[15][14] ;
 wire \core.cpuregs[15][15] ;
 wire \core.cpuregs[15][16] ;
 wire \core.cpuregs[15][17] ;
 wire \core.cpuregs[15][18] ;
 wire \core.cpuregs[15][19] ;
 wire \core.cpuregs[15][1] ;
 wire \core.cpuregs[15][20] ;
 wire \core.cpuregs[15][21] ;
 wire \core.cpuregs[15][22] ;
 wire \core.cpuregs[15][23] ;
 wire \core.cpuregs[15][24] ;
 wire \core.cpuregs[15][25] ;
 wire \core.cpuregs[15][26] ;
 wire \core.cpuregs[15][27] ;
 wire \core.cpuregs[15][28] ;
 wire \core.cpuregs[15][29] ;
 wire \core.cpuregs[15][2] ;
 wire \core.cpuregs[15][30] ;
 wire \core.cpuregs[15][31] ;
 wire \core.cpuregs[15][3] ;
 wire \core.cpuregs[15][4] ;
 wire \core.cpuregs[15][5] ;
 wire \core.cpuregs[15][6] ;
 wire \core.cpuregs[15][7] ;
 wire \core.cpuregs[15][8] ;
 wire \core.cpuregs[15][9] ;
 wire \core.cpuregs[16][0] ;
 wire \core.cpuregs[16][10] ;
 wire \core.cpuregs[16][11] ;
 wire \core.cpuregs[16][12] ;
 wire \core.cpuregs[16][13] ;
 wire \core.cpuregs[16][14] ;
 wire \core.cpuregs[16][15] ;
 wire \core.cpuregs[16][16] ;
 wire \core.cpuregs[16][17] ;
 wire \core.cpuregs[16][18] ;
 wire \core.cpuregs[16][19] ;
 wire \core.cpuregs[16][1] ;
 wire \core.cpuregs[16][20] ;
 wire \core.cpuregs[16][21] ;
 wire \core.cpuregs[16][22] ;
 wire \core.cpuregs[16][23] ;
 wire \core.cpuregs[16][24] ;
 wire \core.cpuregs[16][25] ;
 wire \core.cpuregs[16][26] ;
 wire \core.cpuregs[16][27] ;
 wire \core.cpuregs[16][28] ;
 wire \core.cpuregs[16][29] ;
 wire \core.cpuregs[16][2] ;
 wire \core.cpuregs[16][30] ;
 wire \core.cpuregs[16][31] ;
 wire \core.cpuregs[16][3] ;
 wire \core.cpuregs[16][4] ;
 wire \core.cpuregs[16][5] ;
 wire \core.cpuregs[16][6] ;
 wire \core.cpuregs[16][7] ;
 wire \core.cpuregs[16][8] ;
 wire \core.cpuregs[16][9] ;
 wire \core.cpuregs[17][0] ;
 wire \core.cpuregs[17][10] ;
 wire \core.cpuregs[17][11] ;
 wire \core.cpuregs[17][12] ;
 wire \core.cpuregs[17][13] ;
 wire \core.cpuregs[17][14] ;
 wire \core.cpuregs[17][15] ;
 wire \core.cpuregs[17][16] ;
 wire \core.cpuregs[17][17] ;
 wire \core.cpuregs[17][18] ;
 wire \core.cpuregs[17][19] ;
 wire \core.cpuregs[17][1] ;
 wire \core.cpuregs[17][20] ;
 wire \core.cpuregs[17][21] ;
 wire \core.cpuregs[17][22] ;
 wire \core.cpuregs[17][23] ;
 wire \core.cpuregs[17][24] ;
 wire \core.cpuregs[17][25] ;
 wire \core.cpuregs[17][26] ;
 wire \core.cpuregs[17][27] ;
 wire \core.cpuregs[17][28] ;
 wire \core.cpuregs[17][29] ;
 wire \core.cpuregs[17][2] ;
 wire \core.cpuregs[17][30] ;
 wire \core.cpuregs[17][31] ;
 wire \core.cpuregs[17][3] ;
 wire \core.cpuregs[17][4] ;
 wire \core.cpuregs[17][5] ;
 wire \core.cpuregs[17][6] ;
 wire \core.cpuregs[17][7] ;
 wire \core.cpuregs[17][8] ;
 wire \core.cpuregs[17][9] ;
 wire \core.cpuregs[18][0] ;
 wire \core.cpuregs[18][10] ;
 wire \core.cpuregs[18][11] ;
 wire \core.cpuregs[18][12] ;
 wire \core.cpuregs[18][13] ;
 wire \core.cpuregs[18][14] ;
 wire \core.cpuregs[18][15] ;
 wire \core.cpuregs[18][16] ;
 wire \core.cpuregs[18][17] ;
 wire \core.cpuregs[18][18] ;
 wire \core.cpuregs[18][19] ;
 wire \core.cpuregs[18][1] ;
 wire \core.cpuregs[18][20] ;
 wire \core.cpuregs[18][21] ;
 wire \core.cpuregs[18][22] ;
 wire \core.cpuregs[18][23] ;
 wire \core.cpuregs[18][24] ;
 wire \core.cpuregs[18][25] ;
 wire \core.cpuregs[18][26] ;
 wire \core.cpuregs[18][27] ;
 wire \core.cpuregs[18][28] ;
 wire \core.cpuregs[18][29] ;
 wire \core.cpuregs[18][2] ;
 wire \core.cpuregs[18][30] ;
 wire \core.cpuregs[18][31] ;
 wire \core.cpuregs[18][3] ;
 wire \core.cpuregs[18][4] ;
 wire \core.cpuregs[18][5] ;
 wire \core.cpuregs[18][6] ;
 wire \core.cpuregs[18][7] ;
 wire \core.cpuregs[18][8] ;
 wire \core.cpuregs[18][9] ;
 wire \core.cpuregs[19][0] ;
 wire \core.cpuregs[19][10] ;
 wire \core.cpuregs[19][11] ;
 wire \core.cpuregs[19][12] ;
 wire \core.cpuregs[19][13] ;
 wire \core.cpuregs[19][14] ;
 wire \core.cpuregs[19][15] ;
 wire \core.cpuregs[19][16] ;
 wire \core.cpuregs[19][17] ;
 wire \core.cpuregs[19][18] ;
 wire \core.cpuregs[19][19] ;
 wire \core.cpuregs[19][1] ;
 wire \core.cpuregs[19][20] ;
 wire \core.cpuregs[19][21] ;
 wire \core.cpuregs[19][22] ;
 wire \core.cpuregs[19][23] ;
 wire \core.cpuregs[19][24] ;
 wire \core.cpuregs[19][25] ;
 wire \core.cpuregs[19][26] ;
 wire \core.cpuregs[19][27] ;
 wire \core.cpuregs[19][28] ;
 wire \core.cpuregs[19][29] ;
 wire \core.cpuregs[19][2] ;
 wire \core.cpuregs[19][30] ;
 wire \core.cpuregs[19][31] ;
 wire \core.cpuregs[19][3] ;
 wire \core.cpuregs[19][4] ;
 wire \core.cpuregs[19][5] ;
 wire \core.cpuregs[19][6] ;
 wire \core.cpuregs[19][7] ;
 wire \core.cpuregs[19][8] ;
 wire \core.cpuregs[19][9] ;
 wire \core.cpuregs[1][0] ;
 wire \core.cpuregs[1][10] ;
 wire \core.cpuregs[1][11] ;
 wire \core.cpuregs[1][12] ;
 wire \core.cpuregs[1][13] ;
 wire \core.cpuregs[1][14] ;
 wire \core.cpuregs[1][15] ;
 wire \core.cpuregs[1][16] ;
 wire \core.cpuregs[1][17] ;
 wire \core.cpuregs[1][18] ;
 wire \core.cpuregs[1][19] ;
 wire \core.cpuregs[1][1] ;
 wire \core.cpuregs[1][20] ;
 wire \core.cpuregs[1][21] ;
 wire \core.cpuregs[1][22] ;
 wire \core.cpuregs[1][23] ;
 wire \core.cpuregs[1][24] ;
 wire \core.cpuregs[1][25] ;
 wire \core.cpuregs[1][26] ;
 wire \core.cpuregs[1][27] ;
 wire \core.cpuregs[1][28] ;
 wire \core.cpuregs[1][29] ;
 wire \core.cpuregs[1][2] ;
 wire \core.cpuregs[1][30] ;
 wire \core.cpuregs[1][31] ;
 wire \core.cpuregs[1][3] ;
 wire \core.cpuregs[1][4] ;
 wire \core.cpuregs[1][5] ;
 wire \core.cpuregs[1][6] ;
 wire \core.cpuregs[1][7] ;
 wire \core.cpuregs[1][8] ;
 wire \core.cpuregs[1][9] ;
 wire \core.cpuregs[20][0] ;
 wire \core.cpuregs[20][10] ;
 wire \core.cpuregs[20][11] ;
 wire \core.cpuregs[20][12] ;
 wire \core.cpuregs[20][13] ;
 wire \core.cpuregs[20][14] ;
 wire \core.cpuregs[20][15] ;
 wire \core.cpuregs[20][16] ;
 wire \core.cpuregs[20][17] ;
 wire \core.cpuregs[20][18] ;
 wire \core.cpuregs[20][19] ;
 wire \core.cpuregs[20][1] ;
 wire \core.cpuregs[20][20] ;
 wire \core.cpuregs[20][21] ;
 wire \core.cpuregs[20][22] ;
 wire \core.cpuregs[20][23] ;
 wire \core.cpuregs[20][24] ;
 wire \core.cpuregs[20][25] ;
 wire \core.cpuregs[20][26] ;
 wire \core.cpuregs[20][27] ;
 wire \core.cpuregs[20][28] ;
 wire \core.cpuregs[20][29] ;
 wire \core.cpuregs[20][2] ;
 wire \core.cpuregs[20][30] ;
 wire \core.cpuregs[20][31] ;
 wire \core.cpuregs[20][3] ;
 wire \core.cpuregs[20][4] ;
 wire \core.cpuregs[20][5] ;
 wire \core.cpuregs[20][6] ;
 wire \core.cpuregs[20][7] ;
 wire \core.cpuregs[20][8] ;
 wire \core.cpuregs[20][9] ;
 wire \core.cpuregs[21][0] ;
 wire \core.cpuregs[21][10] ;
 wire \core.cpuregs[21][11] ;
 wire \core.cpuregs[21][12] ;
 wire \core.cpuregs[21][13] ;
 wire \core.cpuregs[21][14] ;
 wire \core.cpuregs[21][15] ;
 wire \core.cpuregs[21][16] ;
 wire \core.cpuregs[21][17] ;
 wire \core.cpuregs[21][18] ;
 wire \core.cpuregs[21][19] ;
 wire \core.cpuregs[21][1] ;
 wire \core.cpuregs[21][20] ;
 wire \core.cpuregs[21][21] ;
 wire \core.cpuregs[21][22] ;
 wire \core.cpuregs[21][23] ;
 wire \core.cpuregs[21][24] ;
 wire \core.cpuregs[21][25] ;
 wire \core.cpuregs[21][26] ;
 wire \core.cpuregs[21][27] ;
 wire \core.cpuregs[21][28] ;
 wire \core.cpuregs[21][29] ;
 wire \core.cpuregs[21][2] ;
 wire \core.cpuregs[21][30] ;
 wire \core.cpuregs[21][31] ;
 wire \core.cpuregs[21][3] ;
 wire \core.cpuregs[21][4] ;
 wire \core.cpuregs[21][5] ;
 wire \core.cpuregs[21][6] ;
 wire \core.cpuregs[21][7] ;
 wire \core.cpuregs[21][8] ;
 wire \core.cpuregs[21][9] ;
 wire \core.cpuregs[22][0] ;
 wire \core.cpuregs[22][10] ;
 wire \core.cpuregs[22][11] ;
 wire \core.cpuregs[22][12] ;
 wire \core.cpuregs[22][13] ;
 wire \core.cpuregs[22][14] ;
 wire \core.cpuregs[22][15] ;
 wire \core.cpuregs[22][16] ;
 wire \core.cpuregs[22][17] ;
 wire \core.cpuregs[22][18] ;
 wire \core.cpuregs[22][19] ;
 wire \core.cpuregs[22][1] ;
 wire \core.cpuregs[22][20] ;
 wire \core.cpuregs[22][21] ;
 wire \core.cpuregs[22][22] ;
 wire \core.cpuregs[22][23] ;
 wire \core.cpuregs[22][24] ;
 wire \core.cpuregs[22][25] ;
 wire \core.cpuregs[22][26] ;
 wire \core.cpuregs[22][27] ;
 wire \core.cpuregs[22][28] ;
 wire \core.cpuregs[22][29] ;
 wire \core.cpuregs[22][2] ;
 wire \core.cpuregs[22][30] ;
 wire \core.cpuregs[22][31] ;
 wire \core.cpuregs[22][3] ;
 wire \core.cpuregs[22][4] ;
 wire \core.cpuregs[22][5] ;
 wire \core.cpuregs[22][6] ;
 wire \core.cpuregs[22][7] ;
 wire \core.cpuregs[22][8] ;
 wire \core.cpuregs[22][9] ;
 wire \core.cpuregs[23][0] ;
 wire \core.cpuregs[23][10] ;
 wire \core.cpuregs[23][11] ;
 wire \core.cpuregs[23][12] ;
 wire \core.cpuregs[23][13] ;
 wire \core.cpuregs[23][14] ;
 wire \core.cpuregs[23][15] ;
 wire \core.cpuregs[23][16] ;
 wire \core.cpuregs[23][17] ;
 wire \core.cpuregs[23][18] ;
 wire \core.cpuregs[23][19] ;
 wire \core.cpuregs[23][1] ;
 wire \core.cpuregs[23][20] ;
 wire \core.cpuregs[23][21] ;
 wire \core.cpuregs[23][22] ;
 wire \core.cpuregs[23][23] ;
 wire \core.cpuregs[23][24] ;
 wire \core.cpuregs[23][25] ;
 wire \core.cpuregs[23][26] ;
 wire \core.cpuregs[23][27] ;
 wire \core.cpuregs[23][28] ;
 wire \core.cpuregs[23][29] ;
 wire \core.cpuregs[23][2] ;
 wire \core.cpuregs[23][30] ;
 wire \core.cpuregs[23][31] ;
 wire \core.cpuregs[23][3] ;
 wire \core.cpuregs[23][4] ;
 wire \core.cpuregs[23][5] ;
 wire \core.cpuregs[23][6] ;
 wire \core.cpuregs[23][7] ;
 wire \core.cpuregs[23][8] ;
 wire \core.cpuregs[23][9] ;
 wire \core.cpuregs[24][0] ;
 wire \core.cpuregs[24][10] ;
 wire \core.cpuregs[24][11] ;
 wire \core.cpuregs[24][12] ;
 wire \core.cpuregs[24][13] ;
 wire \core.cpuregs[24][14] ;
 wire \core.cpuregs[24][15] ;
 wire \core.cpuregs[24][16] ;
 wire \core.cpuregs[24][17] ;
 wire \core.cpuregs[24][18] ;
 wire \core.cpuregs[24][19] ;
 wire \core.cpuregs[24][1] ;
 wire \core.cpuregs[24][20] ;
 wire \core.cpuregs[24][21] ;
 wire \core.cpuregs[24][22] ;
 wire \core.cpuregs[24][23] ;
 wire \core.cpuregs[24][24] ;
 wire \core.cpuregs[24][25] ;
 wire \core.cpuregs[24][26] ;
 wire \core.cpuregs[24][27] ;
 wire \core.cpuregs[24][28] ;
 wire \core.cpuregs[24][29] ;
 wire \core.cpuregs[24][2] ;
 wire \core.cpuregs[24][30] ;
 wire \core.cpuregs[24][31] ;
 wire \core.cpuregs[24][3] ;
 wire \core.cpuregs[24][4] ;
 wire \core.cpuregs[24][5] ;
 wire \core.cpuregs[24][6] ;
 wire \core.cpuregs[24][7] ;
 wire \core.cpuregs[24][8] ;
 wire \core.cpuregs[24][9] ;
 wire \core.cpuregs[25][0] ;
 wire \core.cpuregs[25][10] ;
 wire \core.cpuregs[25][11] ;
 wire \core.cpuregs[25][12] ;
 wire \core.cpuregs[25][13] ;
 wire \core.cpuregs[25][14] ;
 wire \core.cpuregs[25][15] ;
 wire \core.cpuregs[25][16] ;
 wire \core.cpuregs[25][17] ;
 wire \core.cpuregs[25][18] ;
 wire \core.cpuregs[25][19] ;
 wire \core.cpuregs[25][1] ;
 wire \core.cpuregs[25][20] ;
 wire \core.cpuregs[25][21] ;
 wire \core.cpuregs[25][22] ;
 wire \core.cpuregs[25][23] ;
 wire \core.cpuregs[25][24] ;
 wire \core.cpuregs[25][25] ;
 wire \core.cpuregs[25][26] ;
 wire \core.cpuregs[25][27] ;
 wire \core.cpuregs[25][28] ;
 wire \core.cpuregs[25][29] ;
 wire \core.cpuregs[25][2] ;
 wire \core.cpuregs[25][30] ;
 wire \core.cpuregs[25][31] ;
 wire \core.cpuregs[25][3] ;
 wire \core.cpuregs[25][4] ;
 wire \core.cpuregs[25][5] ;
 wire \core.cpuregs[25][6] ;
 wire \core.cpuregs[25][7] ;
 wire \core.cpuregs[25][8] ;
 wire \core.cpuregs[25][9] ;
 wire \core.cpuregs[26][0] ;
 wire \core.cpuregs[26][10] ;
 wire \core.cpuregs[26][11] ;
 wire \core.cpuregs[26][12] ;
 wire \core.cpuregs[26][13] ;
 wire \core.cpuregs[26][14] ;
 wire \core.cpuregs[26][15] ;
 wire \core.cpuregs[26][16] ;
 wire \core.cpuregs[26][17] ;
 wire \core.cpuregs[26][18] ;
 wire \core.cpuregs[26][19] ;
 wire \core.cpuregs[26][1] ;
 wire \core.cpuregs[26][20] ;
 wire \core.cpuregs[26][21] ;
 wire \core.cpuregs[26][22] ;
 wire \core.cpuregs[26][23] ;
 wire \core.cpuregs[26][24] ;
 wire \core.cpuregs[26][25] ;
 wire \core.cpuregs[26][26] ;
 wire \core.cpuregs[26][27] ;
 wire \core.cpuregs[26][28] ;
 wire \core.cpuregs[26][29] ;
 wire \core.cpuregs[26][2] ;
 wire \core.cpuregs[26][30] ;
 wire \core.cpuregs[26][31] ;
 wire \core.cpuregs[26][3] ;
 wire \core.cpuregs[26][4] ;
 wire \core.cpuregs[26][5] ;
 wire \core.cpuregs[26][6] ;
 wire \core.cpuregs[26][7] ;
 wire \core.cpuregs[26][8] ;
 wire \core.cpuregs[26][9] ;
 wire \core.cpuregs[27][0] ;
 wire \core.cpuregs[27][10] ;
 wire \core.cpuregs[27][11] ;
 wire \core.cpuregs[27][12] ;
 wire \core.cpuregs[27][13] ;
 wire \core.cpuregs[27][14] ;
 wire \core.cpuregs[27][15] ;
 wire \core.cpuregs[27][16] ;
 wire \core.cpuregs[27][17] ;
 wire \core.cpuregs[27][18] ;
 wire \core.cpuregs[27][19] ;
 wire \core.cpuregs[27][1] ;
 wire \core.cpuregs[27][20] ;
 wire \core.cpuregs[27][21] ;
 wire \core.cpuregs[27][22] ;
 wire \core.cpuregs[27][23] ;
 wire \core.cpuregs[27][24] ;
 wire \core.cpuregs[27][25] ;
 wire \core.cpuregs[27][26] ;
 wire \core.cpuregs[27][27] ;
 wire \core.cpuregs[27][28] ;
 wire \core.cpuregs[27][29] ;
 wire \core.cpuregs[27][2] ;
 wire \core.cpuregs[27][30] ;
 wire \core.cpuregs[27][31] ;
 wire \core.cpuregs[27][3] ;
 wire \core.cpuregs[27][4] ;
 wire \core.cpuregs[27][5] ;
 wire \core.cpuregs[27][6] ;
 wire \core.cpuregs[27][7] ;
 wire \core.cpuregs[27][8] ;
 wire \core.cpuregs[27][9] ;
 wire \core.cpuregs[28][0] ;
 wire \core.cpuregs[28][10] ;
 wire \core.cpuregs[28][11] ;
 wire \core.cpuregs[28][12] ;
 wire \core.cpuregs[28][13] ;
 wire \core.cpuregs[28][14] ;
 wire \core.cpuregs[28][15] ;
 wire \core.cpuregs[28][16] ;
 wire \core.cpuregs[28][17] ;
 wire \core.cpuregs[28][18] ;
 wire \core.cpuregs[28][19] ;
 wire \core.cpuregs[28][1] ;
 wire \core.cpuregs[28][20] ;
 wire \core.cpuregs[28][21] ;
 wire \core.cpuregs[28][22] ;
 wire \core.cpuregs[28][23] ;
 wire \core.cpuregs[28][24] ;
 wire \core.cpuregs[28][25] ;
 wire \core.cpuregs[28][26] ;
 wire \core.cpuregs[28][27] ;
 wire \core.cpuregs[28][28] ;
 wire \core.cpuregs[28][29] ;
 wire \core.cpuregs[28][2] ;
 wire \core.cpuregs[28][30] ;
 wire \core.cpuregs[28][31] ;
 wire \core.cpuregs[28][3] ;
 wire \core.cpuregs[28][4] ;
 wire \core.cpuregs[28][5] ;
 wire \core.cpuregs[28][6] ;
 wire \core.cpuregs[28][7] ;
 wire \core.cpuregs[28][8] ;
 wire \core.cpuregs[28][9] ;
 wire \core.cpuregs[29][0] ;
 wire \core.cpuregs[29][10] ;
 wire \core.cpuregs[29][11] ;
 wire \core.cpuregs[29][12] ;
 wire \core.cpuregs[29][13] ;
 wire \core.cpuregs[29][14] ;
 wire \core.cpuregs[29][15] ;
 wire \core.cpuregs[29][16] ;
 wire \core.cpuregs[29][17] ;
 wire \core.cpuregs[29][18] ;
 wire \core.cpuregs[29][19] ;
 wire \core.cpuregs[29][1] ;
 wire \core.cpuregs[29][20] ;
 wire \core.cpuregs[29][21] ;
 wire \core.cpuregs[29][22] ;
 wire \core.cpuregs[29][23] ;
 wire \core.cpuregs[29][24] ;
 wire \core.cpuregs[29][25] ;
 wire \core.cpuregs[29][26] ;
 wire \core.cpuregs[29][27] ;
 wire \core.cpuregs[29][28] ;
 wire \core.cpuregs[29][29] ;
 wire \core.cpuregs[29][2] ;
 wire \core.cpuregs[29][30] ;
 wire \core.cpuregs[29][31] ;
 wire \core.cpuregs[29][3] ;
 wire \core.cpuregs[29][4] ;
 wire \core.cpuregs[29][5] ;
 wire \core.cpuregs[29][6] ;
 wire \core.cpuregs[29][7] ;
 wire \core.cpuregs[29][8] ;
 wire \core.cpuregs[29][9] ;
 wire \core.cpuregs[2][0] ;
 wire \core.cpuregs[2][10] ;
 wire \core.cpuregs[2][11] ;
 wire \core.cpuregs[2][12] ;
 wire \core.cpuregs[2][13] ;
 wire \core.cpuregs[2][14] ;
 wire \core.cpuregs[2][15] ;
 wire \core.cpuregs[2][16] ;
 wire \core.cpuregs[2][17] ;
 wire \core.cpuregs[2][18] ;
 wire \core.cpuregs[2][19] ;
 wire \core.cpuregs[2][1] ;
 wire \core.cpuregs[2][20] ;
 wire \core.cpuregs[2][21] ;
 wire \core.cpuregs[2][22] ;
 wire \core.cpuregs[2][23] ;
 wire \core.cpuregs[2][24] ;
 wire \core.cpuregs[2][25] ;
 wire \core.cpuregs[2][26] ;
 wire \core.cpuregs[2][27] ;
 wire \core.cpuregs[2][28] ;
 wire \core.cpuregs[2][29] ;
 wire \core.cpuregs[2][2] ;
 wire \core.cpuregs[2][30] ;
 wire \core.cpuregs[2][31] ;
 wire \core.cpuregs[2][3] ;
 wire \core.cpuregs[2][4] ;
 wire \core.cpuregs[2][5] ;
 wire \core.cpuregs[2][6] ;
 wire \core.cpuregs[2][7] ;
 wire \core.cpuregs[2][8] ;
 wire \core.cpuregs[2][9] ;
 wire \core.cpuregs[30][0] ;
 wire \core.cpuregs[30][10] ;
 wire \core.cpuregs[30][11] ;
 wire \core.cpuregs[30][12] ;
 wire \core.cpuregs[30][13] ;
 wire \core.cpuregs[30][14] ;
 wire \core.cpuregs[30][15] ;
 wire \core.cpuregs[30][16] ;
 wire \core.cpuregs[30][17] ;
 wire \core.cpuregs[30][18] ;
 wire \core.cpuregs[30][19] ;
 wire \core.cpuregs[30][1] ;
 wire \core.cpuregs[30][20] ;
 wire \core.cpuregs[30][21] ;
 wire \core.cpuregs[30][22] ;
 wire \core.cpuregs[30][23] ;
 wire \core.cpuregs[30][24] ;
 wire \core.cpuregs[30][25] ;
 wire \core.cpuregs[30][26] ;
 wire \core.cpuregs[30][27] ;
 wire \core.cpuregs[30][28] ;
 wire \core.cpuregs[30][29] ;
 wire \core.cpuregs[30][2] ;
 wire \core.cpuregs[30][30] ;
 wire \core.cpuregs[30][31] ;
 wire \core.cpuregs[30][3] ;
 wire \core.cpuregs[30][4] ;
 wire \core.cpuregs[30][5] ;
 wire \core.cpuregs[30][6] ;
 wire \core.cpuregs[30][7] ;
 wire \core.cpuregs[30][8] ;
 wire \core.cpuregs[30][9] ;
 wire \core.cpuregs[31][0] ;
 wire \core.cpuregs[31][10] ;
 wire \core.cpuregs[31][11] ;
 wire \core.cpuregs[31][12] ;
 wire \core.cpuregs[31][13] ;
 wire \core.cpuregs[31][14] ;
 wire \core.cpuregs[31][15] ;
 wire \core.cpuregs[31][16] ;
 wire \core.cpuregs[31][17] ;
 wire \core.cpuregs[31][18] ;
 wire \core.cpuregs[31][19] ;
 wire \core.cpuregs[31][1] ;
 wire \core.cpuregs[31][20] ;
 wire \core.cpuregs[31][21] ;
 wire \core.cpuregs[31][22] ;
 wire \core.cpuregs[31][23] ;
 wire \core.cpuregs[31][24] ;
 wire \core.cpuregs[31][25] ;
 wire \core.cpuregs[31][26] ;
 wire \core.cpuregs[31][27] ;
 wire \core.cpuregs[31][28] ;
 wire \core.cpuregs[31][29] ;
 wire \core.cpuregs[31][2] ;
 wire \core.cpuregs[31][30] ;
 wire \core.cpuregs[31][31] ;
 wire \core.cpuregs[31][3] ;
 wire \core.cpuregs[31][4] ;
 wire \core.cpuregs[31][5] ;
 wire \core.cpuregs[31][6] ;
 wire \core.cpuregs[31][7] ;
 wire \core.cpuregs[31][8] ;
 wire \core.cpuregs[31][9] ;
 wire \core.cpuregs[3][0] ;
 wire \core.cpuregs[3][10] ;
 wire \core.cpuregs[3][11] ;
 wire \core.cpuregs[3][12] ;
 wire \core.cpuregs[3][13] ;
 wire \core.cpuregs[3][14] ;
 wire \core.cpuregs[3][15] ;
 wire \core.cpuregs[3][16] ;
 wire \core.cpuregs[3][17] ;
 wire \core.cpuregs[3][18] ;
 wire \core.cpuregs[3][19] ;
 wire \core.cpuregs[3][1] ;
 wire \core.cpuregs[3][20] ;
 wire \core.cpuregs[3][21] ;
 wire \core.cpuregs[3][22] ;
 wire \core.cpuregs[3][23] ;
 wire \core.cpuregs[3][24] ;
 wire \core.cpuregs[3][25] ;
 wire \core.cpuregs[3][26] ;
 wire \core.cpuregs[3][27] ;
 wire \core.cpuregs[3][28] ;
 wire \core.cpuregs[3][29] ;
 wire \core.cpuregs[3][2] ;
 wire \core.cpuregs[3][30] ;
 wire \core.cpuregs[3][31] ;
 wire \core.cpuregs[3][3] ;
 wire \core.cpuregs[3][4] ;
 wire \core.cpuregs[3][5] ;
 wire \core.cpuregs[3][6] ;
 wire \core.cpuregs[3][7] ;
 wire \core.cpuregs[3][8] ;
 wire \core.cpuregs[3][9] ;
 wire \core.cpuregs[4][0] ;
 wire \core.cpuregs[4][10] ;
 wire \core.cpuregs[4][11] ;
 wire \core.cpuregs[4][12] ;
 wire \core.cpuregs[4][13] ;
 wire \core.cpuregs[4][14] ;
 wire \core.cpuregs[4][15] ;
 wire \core.cpuregs[4][16] ;
 wire \core.cpuregs[4][17] ;
 wire \core.cpuregs[4][18] ;
 wire \core.cpuregs[4][19] ;
 wire \core.cpuregs[4][1] ;
 wire \core.cpuregs[4][20] ;
 wire \core.cpuregs[4][21] ;
 wire \core.cpuregs[4][22] ;
 wire \core.cpuregs[4][23] ;
 wire \core.cpuregs[4][24] ;
 wire \core.cpuregs[4][25] ;
 wire \core.cpuregs[4][26] ;
 wire \core.cpuregs[4][27] ;
 wire \core.cpuregs[4][28] ;
 wire \core.cpuregs[4][29] ;
 wire \core.cpuregs[4][2] ;
 wire \core.cpuregs[4][30] ;
 wire \core.cpuregs[4][31] ;
 wire \core.cpuregs[4][3] ;
 wire \core.cpuregs[4][4] ;
 wire \core.cpuregs[4][5] ;
 wire \core.cpuregs[4][6] ;
 wire \core.cpuregs[4][7] ;
 wire \core.cpuregs[4][8] ;
 wire \core.cpuregs[4][9] ;
 wire \core.cpuregs[5][0] ;
 wire \core.cpuregs[5][10] ;
 wire \core.cpuregs[5][11] ;
 wire \core.cpuregs[5][12] ;
 wire \core.cpuregs[5][13] ;
 wire \core.cpuregs[5][14] ;
 wire \core.cpuregs[5][15] ;
 wire \core.cpuregs[5][16] ;
 wire \core.cpuregs[5][17] ;
 wire \core.cpuregs[5][18] ;
 wire \core.cpuregs[5][19] ;
 wire \core.cpuregs[5][1] ;
 wire \core.cpuregs[5][20] ;
 wire \core.cpuregs[5][21] ;
 wire \core.cpuregs[5][22] ;
 wire \core.cpuregs[5][23] ;
 wire \core.cpuregs[5][24] ;
 wire \core.cpuregs[5][25] ;
 wire \core.cpuregs[5][26] ;
 wire \core.cpuregs[5][27] ;
 wire \core.cpuregs[5][28] ;
 wire \core.cpuregs[5][29] ;
 wire \core.cpuregs[5][2] ;
 wire \core.cpuregs[5][30] ;
 wire \core.cpuregs[5][31] ;
 wire \core.cpuregs[5][3] ;
 wire \core.cpuregs[5][4] ;
 wire \core.cpuregs[5][5] ;
 wire \core.cpuregs[5][6] ;
 wire \core.cpuregs[5][7] ;
 wire \core.cpuregs[5][8] ;
 wire \core.cpuregs[5][9] ;
 wire \core.cpuregs[6][0] ;
 wire \core.cpuregs[6][10] ;
 wire \core.cpuregs[6][11] ;
 wire \core.cpuregs[6][12] ;
 wire \core.cpuregs[6][13] ;
 wire \core.cpuregs[6][14] ;
 wire \core.cpuregs[6][15] ;
 wire \core.cpuregs[6][16] ;
 wire \core.cpuregs[6][17] ;
 wire \core.cpuregs[6][18] ;
 wire \core.cpuregs[6][19] ;
 wire \core.cpuregs[6][1] ;
 wire \core.cpuregs[6][20] ;
 wire \core.cpuregs[6][21] ;
 wire \core.cpuregs[6][22] ;
 wire \core.cpuregs[6][23] ;
 wire \core.cpuregs[6][24] ;
 wire \core.cpuregs[6][25] ;
 wire \core.cpuregs[6][26] ;
 wire \core.cpuregs[6][27] ;
 wire \core.cpuregs[6][28] ;
 wire \core.cpuregs[6][29] ;
 wire \core.cpuregs[6][2] ;
 wire \core.cpuregs[6][30] ;
 wire \core.cpuregs[6][31] ;
 wire \core.cpuregs[6][3] ;
 wire \core.cpuregs[6][4] ;
 wire \core.cpuregs[6][5] ;
 wire \core.cpuregs[6][6] ;
 wire \core.cpuregs[6][7] ;
 wire \core.cpuregs[6][8] ;
 wire \core.cpuregs[6][9] ;
 wire \core.cpuregs[7][0] ;
 wire \core.cpuregs[7][10] ;
 wire \core.cpuregs[7][11] ;
 wire \core.cpuregs[7][12] ;
 wire \core.cpuregs[7][13] ;
 wire \core.cpuregs[7][14] ;
 wire \core.cpuregs[7][15] ;
 wire \core.cpuregs[7][16] ;
 wire \core.cpuregs[7][17] ;
 wire \core.cpuregs[7][18] ;
 wire \core.cpuregs[7][19] ;
 wire \core.cpuregs[7][1] ;
 wire \core.cpuregs[7][20] ;
 wire \core.cpuregs[7][21] ;
 wire \core.cpuregs[7][22] ;
 wire \core.cpuregs[7][23] ;
 wire \core.cpuregs[7][24] ;
 wire \core.cpuregs[7][25] ;
 wire \core.cpuregs[7][26] ;
 wire \core.cpuregs[7][27] ;
 wire \core.cpuregs[7][28] ;
 wire \core.cpuregs[7][29] ;
 wire \core.cpuregs[7][2] ;
 wire \core.cpuregs[7][30] ;
 wire \core.cpuregs[7][31] ;
 wire \core.cpuregs[7][3] ;
 wire \core.cpuregs[7][4] ;
 wire \core.cpuregs[7][5] ;
 wire \core.cpuregs[7][6] ;
 wire \core.cpuregs[7][7] ;
 wire \core.cpuregs[7][8] ;
 wire \core.cpuregs[7][9] ;
 wire \core.cpuregs[8][0] ;
 wire \core.cpuregs[8][10] ;
 wire \core.cpuregs[8][11] ;
 wire \core.cpuregs[8][12] ;
 wire \core.cpuregs[8][13] ;
 wire \core.cpuregs[8][14] ;
 wire \core.cpuregs[8][15] ;
 wire \core.cpuregs[8][16] ;
 wire \core.cpuregs[8][17] ;
 wire \core.cpuregs[8][18] ;
 wire \core.cpuregs[8][19] ;
 wire \core.cpuregs[8][1] ;
 wire \core.cpuregs[8][20] ;
 wire \core.cpuregs[8][21] ;
 wire \core.cpuregs[8][22] ;
 wire \core.cpuregs[8][23] ;
 wire \core.cpuregs[8][24] ;
 wire \core.cpuregs[8][25] ;
 wire \core.cpuregs[8][26] ;
 wire \core.cpuregs[8][27] ;
 wire \core.cpuregs[8][28] ;
 wire \core.cpuregs[8][29] ;
 wire \core.cpuregs[8][2] ;
 wire \core.cpuregs[8][30] ;
 wire \core.cpuregs[8][31] ;
 wire \core.cpuregs[8][3] ;
 wire \core.cpuregs[8][4] ;
 wire \core.cpuregs[8][5] ;
 wire \core.cpuregs[8][6] ;
 wire \core.cpuregs[8][7] ;
 wire \core.cpuregs[8][8] ;
 wire \core.cpuregs[8][9] ;
 wire \core.cpuregs[9][0] ;
 wire \core.cpuregs[9][10] ;
 wire \core.cpuregs[9][11] ;
 wire \core.cpuregs[9][12] ;
 wire \core.cpuregs[9][13] ;
 wire \core.cpuregs[9][14] ;
 wire \core.cpuregs[9][15] ;
 wire \core.cpuregs[9][16] ;
 wire \core.cpuregs[9][17] ;
 wire \core.cpuregs[9][18] ;
 wire \core.cpuregs[9][19] ;
 wire \core.cpuregs[9][1] ;
 wire \core.cpuregs[9][20] ;
 wire \core.cpuregs[9][21] ;
 wire \core.cpuregs[9][22] ;
 wire \core.cpuregs[9][23] ;
 wire \core.cpuregs[9][24] ;
 wire \core.cpuregs[9][25] ;
 wire \core.cpuregs[9][26] ;
 wire \core.cpuregs[9][27] ;
 wire \core.cpuregs[9][28] ;
 wire \core.cpuregs[9][29] ;
 wire \core.cpuregs[9][2] ;
 wire \core.cpuregs[9][30] ;
 wire \core.cpuregs[9][31] ;
 wire \core.cpuregs[9][3] ;
 wire \core.cpuregs[9][4] ;
 wire \core.cpuregs[9][5] ;
 wire \core.cpuregs[9][6] ;
 wire \core.cpuregs[9][7] ;
 wire \core.cpuregs[9][8] ;
 wire \core.cpuregs[9][9] ;
 wire \core.decoded_imm[0] ;
 wire \core.decoded_imm[10] ;
 wire \core.decoded_imm[11] ;
 wire \core.decoded_imm[12] ;
 wire \core.decoded_imm[13] ;
 wire \core.decoded_imm[14] ;
 wire \core.decoded_imm[15] ;
 wire \core.decoded_imm[16] ;
 wire \core.decoded_imm[17] ;
 wire \core.decoded_imm[18] ;
 wire \core.decoded_imm[19] ;
 wire \core.decoded_imm[1] ;
 wire \core.decoded_imm[20] ;
 wire \core.decoded_imm[21] ;
 wire \core.decoded_imm[22] ;
 wire \core.decoded_imm[23] ;
 wire \core.decoded_imm[24] ;
 wire \core.decoded_imm[25] ;
 wire \core.decoded_imm[26] ;
 wire \core.decoded_imm[27] ;
 wire \core.decoded_imm[28] ;
 wire \core.decoded_imm[29] ;
 wire \core.decoded_imm[2] ;
 wire \core.decoded_imm[30] ;
 wire \core.decoded_imm[31] ;
 wire \core.decoded_imm[3] ;
 wire \core.decoded_imm[4] ;
 wire \core.decoded_imm[5] ;
 wire \core.decoded_imm[6] ;
 wire \core.decoded_imm[7] ;
 wire \core.decoded_imm[8] ;
 wire \core.decoded_imm[9] ;
 wire \core.decoded_imm_j[10] ;
 wire \core.decoded_imm_j[11] ;
 wire \core.decoded_imm_j[12] ;
 wire \core.decoded_imm_j[13] ;
 wire \core.decoded_imm_j[14] ;
 wire \core.decoded_imm_j[15] ;
 wire \core.decoded_imm_j[16] ;
 wire \core.decoded_imm_j[17] ;
 wire \core.decoded_imm_j[18] ;
 wire \core.decoded_imm_j[19] ;
 wire \core.decoded_imm_j[1] ;
 wire \core.decoded_imm_j[20] ;
 wire \core.decoded_imm_j[2] ;
 wire \core.decoded_imm_j[3] ;
 wire \core.decoded_imm_j[4] ;
 wire \core.decoded_imm_j[5] ;
 wire \core.decoded_imm_j[6] ;
 wire \core.decoded_imm_j[7] ;
 wire \core.decoded_imm_j[8] ;
 wire \core.decoded_imm_j[9] ;
 wire \core.decoded_rd[0] ;
 wire \core.decoded_rd[1] ;
 wire \core.decoded_rd[2] ;
 wire \core.decoded_rd[3] ;
 wire \core.decoded_rd[4] ;
 wire \core.decoder_pseudo_trigger ;
 wire \core.decoder_trigger ;
 wire \core.instr_add ;
 wire \core.instr_addi ;
 wire \core.instr_and ;
 wire \core.instr_andi ;
 wire \core.instr_auipc ;
 wire \core.instr_beq ;
 wire \core.instr_bge ;
 wire \core.instr_bgeu ;
 wire \core.instr_blt ;
 wire \core.instr_bltu ;
 wire \core.instr_bne ;
 wire \core.instr_fence ;
 wire \core.instr_jal ;
 wire \core.instr_jalr ;
 wire \core.instr_lb ;
 wire \core.instr_lbu ;
 wire \core.instr_lh ;
 wire \core.instr_lhu ;
 wire \core.instr_lui ;
 wire \core.instr_lw ;
 wire \core.instr_or ;
 wire \core.instr_ori ;
 wire \core.instr_rdcycle ;
 wire \core.instr_rdcycleh ;
 wire \core.instr_rdinstr ;
 wire \core.instr_rdinstrh ;
 wire \core.instr_sb ;
 wire \core.instr_sh ;
 wire \core.instr_sll ;
 wire \core.instr_slli ;
 wire \core.instr_slt ;
 wire \core.instr_slti ;
 wire \core.instr_sltiu ;
 wire \core.instr_sltu ;
 wire \core.instr_sra ;
 wire \core.instr_srai ;
 wire \core.instr_srl ;
 wire \core.instr_srli ;
 wire \core.instr_sub ;
 wire \core.instr_sw ;
 wire \core.instr_xor ;
 wire \core.instr_xori ;
 wire \core.is_alu_reg_imm ;
 wire \core.is_alu_reg_reg ;
 wire \core.is_beq_bne_blt_bge_bltu_bgeu ;
 wire \core.is_compare ;
 wire \core.is_jalr_addi_slti_sltiu_xori_ori_andi ;
 wire \core.is_lb_lh_lw_lbu_lhu ;
 wire \core.is_lui_auipc_jal ;
 wire \core.is_sb_sh_sw ;
 wire \core.is_sll_srl_sra ;
 wire \core.is_slli_srli_srai ;
 wire \core.is_slti_blt_slt ;
 wire \core.is_sltiu_bltu_sltu ;
 wire \core.latched_branch ;
 wire \core.latched_is_lb ;
 wire \core.latched_is_lh ;
 wire \core.latched_rd[0] ;
 wire \core.latched_rd[1] ;
 wire \core.latched_rd[2] ;
 wire \core.latched_rd[3] ;
 wire \core.latched_rd[4] ;
 wire \core.latched_stalu ;
 wire \core.latched_store ;
 wire \core.mem_do_prefetch ;
 wire \core.mem_do_rdata ;
 wire \core.mem_do_rinst ;
 wire \core.mem_do_wdata ;
 wire \core.mem_la_wdata[0] ;
 wire \core.mem_la_wdata[1] ;
 wire \core.mem_la_wdata[2] ;
 wire \core.mem_la_wdata[3] ;
 wire \core.mem_la_wdata[4] ;
 wire \core.mem_la_wdata[5] ;
 wire \core.mem_la_wdata[6] ;
 wire \core.mem_la_wdata[7] ;
 wire \core.mem_rdata_q[0] ;
 wire \core.mem_rdata_q[10] ;
 wire \core.mem_rdata_q[11] ;
 wire \core.mem_rdata_q[12] ;
 wire \core.mem_rdata_q[13] ;
 wire \core.mem_rdata_q[14] ;
 wire \core.mem_rdata_q[15] ;
 wire \core.mem_rdata_q[16] ;
 wire \core.mem_rdata_q[17] ;
 wire \core.mem_rdata_q[18] ;
 wire \core.mem_rdata_q[19] ;
 wire \core.mem_rdata_q[1] ;
 wire \core.mem_rdata_q[20] ;
 wire \core.mem_rdata_q[21] ;
 wire \core.mem_rdata_q[22] ;
 wire \core.mem_rdata_q[23] ;
 wire \core.mem_rdata_q[24] ;
 wire \core.mem_rdata_q[25] ;
 wire \core.mem_rdata_q[26] ;
 wire \core.mem_rdata_q[27] ;
 wire \core.mem_rdata_q[28] ;
 wire \core.mem_rdata_q[29] ;
 wire \core.mem_rdata_q[2] ;
 wire \core.mem_rdata_q[30] ;
 wire \core.mem_rdata_q[31] ;
 wire \core.mem_rdata_q[3] ;
 wire \core.mem_rdata_q[4] ;
 wire \core.mem_rdata_q[5] ;
 wire \core.mem_rdata_q[6] ;
 wire \core.mem_rdata_q[7] ;
 wire \core.mem_rdata_q[8] ;
 wire \core.mem_rdata_q[9] ;
 wire \core.mem_state[0] ;
 wire \core.mem_state[1] ;
 wire \core.mem_wordsize[0] ;
 wire \core.mem_wordsize[1] ;
 wire \core.mem_wordsize[2] ;
 wire \core.pcpi_rs1[0] ;
 wire \core.pcpi_rs1[10] ;
 wire \core.pcpi_rs1[11] ;
 wire \core.pcpi_rs1[12] ;
 wire \core.pcpi_rs1[13] ;
 wire \core.pcpi_rs1[14] ;
 wire \core.pcpi_rs1[15] ;
 wire \core.pcpi_rs1[16] ;
 wire \core.pcpi_rs1[17] ;
 wire \core.pcpi_rs1[18] ;
 wire \core.pcpi_rs1[19] ;
 wire \core.pcpi_rs1[1] ;
 wire \core.pcpi_rs1[20] ;
 wire \core.pcpi_rs1[21] ;
 wire \core.pcpi_rs1[22] ;
 wire \core.pcpi_rs1[23] ;
 wire \core.pcpi_rs1[24] ;
 wire \core.pcpi_rs1[25] ;
 wire \core.pcpi_rs1[26] ;
 wire \core.pcpi_rs1[27] ;
 wire \core.pcpi_rs1[28] ;
 wire \core.pcpi_rs1[29] ;
 wire \core.pcpi_rs1[2] ;
 wire \core.pcpi_rs1[30] ;
 wire \core.pcpi_rs1[31] ;
 wire \core.pcpi_rs1[3] ;
 wire \core.pcpi_rs1[4] ;
 wire \core.pcpi_rs1[5] ;
 wire \core.pcpi_rs1[6] ;
 wire \core.pcpi_rs1[7] ;
 wire \core.pcpi_rs1[8] ;
 wire \core.pcpi_rs1[9] ;
 wire \core.pcpi_rs2[10] ;
 wire \core.pcpi_rs2[11] ;
 wire \core.pcpi_rs2[12] ;
 wire \core.pcpi_rs2[13] ;
 wire \core.pcpi_rs2[14] ;
 wire \core.pcpi_rs2[15] ;
 wire \core.pcpi_rs2[16] ;
 wire \core.pcpi_rs2[17] ;
 wire \core.pcpi_rs2[18] ;
 wire \core.pcpi_rs2[19] ;
 wire \core.pcpi_rs2[20] ;
 wire \core.pcpi_rs2[21] ;
 wire \core.pcpi_rs2[22] ;
 wire \core.pcpi_rs2[23] ;
 wire \core.pcpi_rs2[24] ;
 wire \core.pcpi_rs2[25] ;
 wire \core.pcpi_rs2[26] ;
 wire \core.pcpi_rs2[27] ;
 wire \core.pcpi_rs2[28] ;
 wire \core.pcpi_rs2[29] ;
 wire \core.pcpi_rs2[30] ;
 wire \core.pcpi_rs2[31] ;
 wire \core.pcpi_rs2[8] ;
 wire \core.pcpi_rs2[9] ;
 wire \core.reg_next_pc[10] ;
 wire \core.reg_next_pc[11] ;
 wire \core.reg_next_pc[12] ;
 wire \core.reg_next_pc[13] ;
 wire \core.reg_next_pc[14] ;
 wire \core.reg_next_pc[15] ;
 wire \core.reg_next_pc[16] ;
 wire \core.reg_next_pc[17] ;
 wire \core.reg_next_pc[18] ;
 wire \core.reg_next_pc[19] ;
 wire \core.reg_next_pc[1] ;
 wire \core.reg_next_pc[20] ;
 wire \core.reg_next_pc[21] ;
 wire \core.reg_next_pc[22] ;
 wire \core.reg_next_pc[23] ;
 wire \core.reg_next_pc[24] ;
 wire \core.reg_next_pc[25] ;
 wire \core.reg_next_pc[26] ;
 wire \core.reg_next_pc[27] ;
 wire \core.reg_next_pc[28] ;
 wire \core.reg_next_pc[29] ;
 wire \core.reg_next_pc[2] ;
 wire \core.reg_next_pc[30] ;
 wire \core.reg_next_pc[31] ;
 wire \core.reg_next_pc[3] ;
 wire \core.reg_next_pc[4] ;
 wire \core.reg_next_pc[5] ;
 wire \core.reg_next_pc[6] ;
 wire \core.reg_next_pc[7] ;
 wire \core.reg_next_pc[8] ;
 wire \core.reg_next_pc[9] ;
 wire \core.reg_out[0] ;
 wire \core.reg_out[10] ;
 wire \core.reg_out[11] ;
 wire \core.reg_out[12] ;
 wire \core.reg_out[13] ;
 wire \core.reg_out[14] ;
 wire \core.reg_out[15] ;
 wire \core.reg_out[16] ;
 wire \core.reg_out[17] ;
 wire \core.reg_out[18] ;
 wire \core.reg_out[19] ;
 wire \core.reg_out[1] ;
 wire \core.reg_out[20] ;
 wire \core.reg_out[21] ;
 wire \core.reg_out[22] ;
 wire \core.reg_out[23] ;
 wire \core.reg_out[24] ;
 wire \core.reg_out[25] ;
 wire \core.reg_out[26] ;
 wire \core.reg_out[27] ;
 wire \core.reg_out[28] ;
 wire \core.reg_out[29] ;
 wire \core.reg_out[2] ;
 wire \core.reg_out[30] ;
 wire \core.reg_out[31] ;
 wire \core.reg_out[3] ;
 wire \core.reg_out[4] ;
 wire \core.reg_out[5] ;
 wire \core.reg_out[6] ;
 wire \core.reg_out[7] ;
 wire \core.reg_out[8] ;
 wire \core.reg_out[9] ;
 wire \core.reg_pc[10] ;
 wire \core.reg_pc[11] ;
 wire \core.reg_pc[12] ;
 wire \core.reg_pc[13] ;
 wire \core.reg_pc[14] ;
 wire \core.reg_pc[15] ;
 wire \core.reg_pc[16] ;
 wire \core.reg_pc[17] ;
 wire \core.reg_pc[18] ;
 wire \core.reg_pc[19] ;
 wire \core.reg_pc[1] ;
 wire \core.reg_pc[20] ;
 wire \core.reg_pc[21] ;
 wire \core.reg_pc[22] ;
 wire \core.reg_pc[23] ;
 wire \core.reg_pc[24] ;
 wire \core.reg_pc[25] ;
 wire \core.reg_pc[26] ;
 wire \core.reg_pc[27] ;
 wire \core.reg_pc[28] ;
 wire \core.reg_pc[29] ;
 wire \core.reg_pc[2] ;
 wire \core.reg_pc[30] ;
 wire \core.reg_pc[31] ;
 wire \core.reg_pc[3] ;
 wire \core.reg_pc[4] ;
 wire \core.reg_pc[5] ;
 wire \core.reg_pc[6] ;
 wire \core.reg_pc[7] ;
 wire \core.reg_pc[8] ;
 wire \core.reg_pc[9] ;
 wire \core.reg_sh[0] ;
 wire \core.reg_sh[1] ;
 wire \core.reg_sh[2] ;
 wire \core.reg_sh[3] ;
 wire \core.reg_sh[4] ;
 wire net107;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;

 sky130_fd_sc_hd__or3_1 _10452_ (.A(\core.instr_sltu ),
    .B(\core.instr_bltu ),
    .C(\core.instr_sltiu ),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _10453_ (.A(_04362_),
    .X(_00033_));
 sky130_fd_sc_hd__or3_1 _10454_ (.A(\core.instr_slt ),
    .B(\core.instr_blt ),
    .C(\core.instr_slti ),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _10455_ (.A(_04363_),
    .X(_00032_));
 sky130_fd_sc_hd__nor2_1 _10456_ (.A(\core.instr_auipc ),
    .B(\core.instr_lui ),
    .Y(_04364_));
 sky130_fd_sc_hd__inv_2 _10457_ (.A(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__nor2_2 _10458_ (.A(\core.instr_jal ),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__inv_2 _10459_ (.A(_04366_),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _10460_ (.A(\core.mem_do_prefetch ),
    .Y(_04367_));
 sky130_fd_sc_hd__inv_2 _10461_ (.A(\core.mem_do_rinst ),
    .Y(_04368_));
 sky130_fd_sc_hd__inv_2 _10462_ (.A(\core.mem_do_rdata ),
    .Y(_04369_));
 sky130_fd_sc_hd__inv_2 _10463_ (.A(\core.mem_do_wdata ),
    .Y(_04370_));
 sky130_fd_sc_hd__nor2_2 _10464_ (.A(\core.mem_state[1] ),
    .B(\core.mem_state[0] ),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _10465_ (.A(net66),
    .B(net33),
    .Y(_04372_));
 sky130_fd_sc_hd__a311o_1 _10466_ (.A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .B1(_04371_),
    .C1(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__inv_2 _10467_ (.A(\core.mem_state[1] ),
    .Y(_04374_));
 sky130_fd_sc_hd__inv_2 _10468_ (.A(\core.mem_state[0] ),
    .Y(_04375_));
 sky130_fd_sc_hd__or3_1 _10469_ (.A(_04368_),
    .B(_04374_),
    .C(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(_04373_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__and2_1 _10471_ (.A(_04377_),
    .B(net34),
    .X(_04378_));
 sky130_fd_sc_hd__nor2_1 _10472_ (.A(_04367_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__inv_2 _10473_ (.A(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_1 _10474_ (.A(_04380_),
    .B(_04370_),
    .Y(_04381_));
 sky130_fd_sc_hd__nand2_1 _10475_ (.A(net34),
    .B(\core.cpu_state[5] ),
    .Y(_04382_));
 sky130_fd_sc_hd__inv_2 _10476_ (.A(\core.instr_sb ),
    .Y(_04383_));
 sky130_fd_sc_hd__inv_2 _10477_ (.A(\core.instr_sh ),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_1 _10478_ (.A(_04383_),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__or3_1 _10479_ (.A(\core.instr_sw ),
    .B(_04382_),
    .C(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_2 _10480_ (.A(net34),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_2 _10481_ (.A(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__and3_1 _10482_ (.A(_04380_),
    .B(\core.mem_do_wdata ),
    .C(\core.cpu_state[5] ),
    .X(_04389_));
 sky130_fd_sc_hd__a2bb2o_1 _10483_ (.A1_N(_04381_),
    .A2_N(_04386_),
    .B1(_04388_),
    .B2(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_2 _10484_ (.A(\core.cpu_state[1] ),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_2 _10485_ (.A(\core.cpu_state[6] ),
    .X(_04392_));
 sky130_fd_sc_hd__nor2_2 _10486_ (.A(_04391_),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__inv_2 _10487_ (.A(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nor2_2 _10488_ (.A(\core.cpu_state[6] ),
    .B(\core.cpu_state[5] ),
    .Y(_04395_));
 sky130_fd_sc_hd__inv_2 _10489_ (.A(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10490_ (.A(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__nand2_1 _10491_ (.A(_04379_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__inv_2 _10492_ (.A(_04392_),
    .Y(_04399_));
 sky130_fd_sc_hd__or3_4 _10493_ (.A(_04369_),
    .B(_04399_),
    .C(_04379_),
    .X(_04400_));
 sky130_fd_sc_hd__o2111a_1 _10494_ (.A1(\core.cpu_state[5] ),
    .A2(_04394_),
    .B1(_04388_),
    .C1(_04398_),
    .D1(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__nor2_1 _10495_ (.A(\core.instr_lb ),
    .B(\core.instr_lbu ),
    .Y(_04402_));
 sky130_fd_sc_hd__inv_2 _10496_ (.A(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__or2_1 _10497_ (.A(\core.instr_lh ),
    .B(\core.instr_lhu ),
    .X(_04404_));
 sky130_fd_sc_hd__or2_1 _10498_ (.A(_04403_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__nand2_1 _10499_ (.A(_04387_),
    .B(_04392_),
    .Y(_04406_));
 sky130_fd_sc_hd__or3_2 _10500_ (.A(\core.mem_do_rdata ),
    .B(_04406_),
    .C(_04379_),
    .X(_04407_));
 sky130_fd_sc_hd__or3_1 _10501_ (.A(\core.instr_lw ),
    .B(_04405_),
    .C(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__nand3b_1 _10502_ (.A_N(_04390_),
    .B(_04401_),
    .C(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__clkbuf_2 _10503_ (.A(\core.mem_wordsize[1] ),
    .X(_04410_));
 sky130_fd_sc_hd__clkbuf_2 _10504_ (.A(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__or3_1 _10505_ (.A(_04383_),
    .B(_04382_),
    .C(_04381_),
    .X(_04412_));
 sky130_fd_sc_hd__o21ai_1 _10506_ (.A1(_04407_),
    .A2(_04402_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a21o_1 _10507_ (.A1(_04409_),
    .A2(_04411_),
    .B1(_04413_),
    .X(_00018_));
 sky130_fd_sc_hd__nor2_1 _10508_ (.A(\core.instr_slt ),
    .B(\core.instr_sltu ),
    .Y(_04414_));
 sky130_fd_sc_hd__or3b_1 _10509_ (.A(_04385_),
    .B(_04403_),
    .C_N(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__or4_1 _10510_ (.A(\core.instr_srl ),
    .B(\core.instr_or ),
    .C(\core.instr_and ),
    .D(\core.instr_blt ),
    .X(_04416_));
 sky130_fd_sc_hd__or4_1 _10511_ (.A(\core.instr_addi ),
    .B(\core.instr_xori ),
    .C(\core.instr_andi ),
    .D(\core.instr_sub ),
    .X(_04417_));
 sky130_fd_sc_hd__or3_1 _10512_ (.A(_04415_),
    .B(_04416_),
    .C(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__or4_1 _10513_ (.A(\core.instr_sll ),
    .B(\core.instr_add ),
    .C(\core.instr_ori ),
    .D(\core.instr_sltiu ),
    .X(_04419_));
 sky130_fd_sc_hd__or4_1 _10514_ (.A(\core.instr_bltu ),
    .B(\core.instr_fence ),
    .C(\core.instr_sra ),
    .D(\core.instr_xor ),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _10515_ (.A(\core.instr_rdcycle ),
    .B(\core.instr_srai ),
    .Y(_04421_));
 sky130_fd_sc_hd__inv_2 _10516_ (.A(\core.instr_slti ),
    .Y(_04422_));
 sky130_fd_sc_hd__inv_2 _10517_ (.A(\core.instr_beq ),
    .Y(_04423_));
 sky130_fd_sc_hd__and3_1 _10518_ (.A(_04421_),
    .B(_04422_),
    .C(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__inv_2 _10519_ (.A(\core.instr_jalr ),
    .Y(_04425_));
 sky130_fd_sc_hd__inv_2 _10520_ (.A(\core.instr_lh ),
    .Y(_04426_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(\core.instr_srli ),
    .B(\core.instr_slli ),
    .Y(_04427_));
 sky130_fd_sc_hd__and4_1 _10522_ (.A(_04424_),
    .B(_04425_),
    .C(_04426_),
    .D(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__or3b_1 _10523_ (.A(_04419_),
    .B(_04420_),
    .C_N(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__nor2_1 _10524_ (.A(_04418_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__or3_2 _10525_ (.A(\core.instr_rdinstr ),
    .B(\core.instr_rdinstrh ),
    .C(\core.instr_rdcycleh ),
    .X(_04431_));
 sky130_fd_sc_hd__inv_2 _10526_ (.A(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nor3_1 _10527_ (.A(\core.instr_lhu ),
    .B(\core.instr_lw ),
    .C(\core.instr_sw ),
    .Y(_04433_));
 sky130_fd_sc_hd__inv_2 _10528_ (.A(\core.instr_bgeu ),
    .Y(_04434_));
 sky130_fd_sc_hd__inv_2 _10529_ (.A(\core.instr_bge ),
    .Y(_04435_));
 sky130_fd_sc_hd__inv_2 _10530_ (.A(\core.instr_bne ),
    .Y(_04436_));
 sky130_fd_sc_hd__and3_1 _10531_ (.A(_04434_),
    .B(_04435_),
    .C(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__and4_1 _10532_ (.A(_04432_),
    .B(_04366_),
    .C(_04433_),
    .D(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__inv_2 _10533_ (.A(\core.cpu_state[2] ),
    .Y(_04439_));
 sky130_fd_sc_hd__clkbuf_2 _10534_ (.A(\core.mem_wordsize[2] ),
    .X(_04440_));
 sky130_fd_sc_hd__clkbuf_2 _10535_ (.A(\core.pcpi_rs1[0] ),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_2 _10536_ (.A(\core.pcpi_rs1[1] ),
    .X(_04442_));
 sky130_fd_sc_hd__nor2_1 _10537_ (.A(_04441_),
    .B(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__inv_2 _10538_ (.A(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__a22o_1 _10539_ (.A1(_04440_),
    .A2(_04441_),
    .B1(_04444_),
    .B2(\core.mem_wordsize[0] ),
    .X(_04445_));
 sky130_fd_sc_hd__o21a_1 _10540_ (.A1(\core.mem_do_rdata ),
    .A2(\core.mem_do_wdata ),
    .B1(_04387_),
    .X(_04446_));
 sky130_fd_sc_hd__and3_1 _10541_ (.A(\core.mem_do_rinst ),
    .B(\core.reg_pc[1] ),
    .C(net34),
    .X(_04447_));
 sky130_fd_sc_hd__a21oi_4 _10542_ (.A1(_04445_),
    .A2(_04446_),
    .B1(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand2_1 _10543_ (.A(_04448_),
    .B(_04387_),
    .Y(_04449_));
 sky130_fd_sc_hd__nor2_1 _10544_ (.A(_04439_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__buf_1 _10545_ (.A(_04387_),
    .X(_04451_));
 sky130_fd_sc_hd__nand2_1 _10546_ (.A(_04451_),
    .B(\core.cpu_state[0] ),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_4 _10547_ (.A(_04448_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__a31o_1 _10548_ (.A1(_04430_),
    .A2(_04438_),
    .A3(_04450_),
    .B1(_04453_),
    .X(_00010_));
 sky130_fd_sc_hd__or3b_1 _10549_ (.A(_04382_),
    .B(_04381_),
    .C_N(\core.instr_sw ),
    .X(_04454_));
 sky130_fd_sc_hd__inv_4 _10550_ (.A(_04407_),
    .Y(_04455_));
 sky130_fd_sc_hd__nand2_1 _10551_ (.A(_04455_),
    .B(\core.instr_lw ),
    .Y(_04456_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(\core.cpu_state[1] ),
    .B(net34),
    .Y(_04457_));
 sky130_fd_sc_hd__and3_1 _10553_ (.A(_04454_),
    .B(_04456_),
    .C(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__a21bo_1 _10554_ (.A1(_04409_),
    .A2(net108),
    .B1_N(_04458_),
    .X(_00017_));
 sky130_fd_sc_hd__clkbuf_2 _10555_ (.A(_04392_),
    .X(_04459_));
 sky130_fd_sc_hd__inv_2 _10556_ (.A(_04449_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _10557_ (.A(_04378_),
    .B(_04367_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(_04430_),
    .B(_04438_),
    .Y(_04462_));
 sky130_fd_sc_hd__and3_1 _10559_ (.A(_04462_),
    .B(\core.is_lb_lh_lw_lbu_lhu ),
    .C(_04450_),
    .X(_04463_));
 sky130_fd_sc_hd__a31o_1 _10560_ (.A1(_04459_),
    .A2(_04460_),
    .A3(_04461_),
    .B1(_04463_),
    .X(_00016_));
 sky130_fd_sc_hd__nand2_1 _10561_ (.A(_04462_),
    .B(\core.is_lb_lh_lw_lbu_lhu ),
    .Y(_04464_));
 sky130_fd_sc_hd__nor2_1 _10562_ (.A(\core.instr_rdcycle ),
    .B(_04431_),
    .Y(_04465_));
 sky130_fd_sc_hd__buf_1 _10563_ (.A(\core.cpu_state[2] ),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_2 _10564_ (.A(\core.is_sb_sh_sw ),
    .X(_04467_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10565_ (.A(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__and3_1 _10566_ (.A(_04465_),
    .B(_04466_),
    .C(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__and3_1 _10567_ (.A(_04464_),
    .B(_04460_),
    .C(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__inv_2 _10568_ (.A(\core.is_slli_srli_srai ),
    .Y(_04471_));
 sky130_fd_sc_hd__and2_1 _10569_ (.A(_04462_),
    .B(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_2 _10570_ (.A(\core.is_lui_auipc_jal ),
    .B(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .Y(_04473_));
 sky130_fd_sc_hd__clkbuf_2 _10571_ (.A(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_04472_),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__inv_2 _10573_ (.A(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__a32o_1 _10574_ (.A1(\core.cpu_state[5] ),
    .A2(_04460_),
    .A3(_04461_),
    .B1(_04470_),
    .B2(_04476_),
    .X(_00015_));
 sky130_fd_sc_hd__inv_2 _10575_ (.A(\core.is_sll_srl_sra ),
    .Y(_04477_));
 sky130_fd_sc_hd__inv_2 _10576_ (.A(_04465_),
    .Y(_04478_));
 sky130_fd_sc_hd__nor2_1 _10577_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__or2_1 _10578_ (.A(\core.reg_sh[3] ),
    .B(\core.reg_sh[2] ),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_1 _10579_ (.A(\core.reg_sh[4] ),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__nor2_1 _10580_ (.A(\core.reg_sh[0] ),
    .B(\core.reg_sh[1] ),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_1 _10581_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_04483_),
    .B(\core.cpu_state[4] ),
    .Y(_04484_));
 sky130_fd_sc_hd__buf_1 _10583_ (.A(\core.is_slli_srli_srai ),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_04466_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__a21oi_1 _10585_ (.A1(_04484_),
    .A2(_04486_),
    .B1(_04449_),
    .Y(_04487_));
 sky130_fd_sc_hd__a41o_1 _10586_ (.A1(_04476_),
    .A2(_04450_),
    .A3(_04464_),
    .A4(_04479_),
    .B1(_04487_),
    .X(_00014_));
 sky130_fd_sc_hd__clkbuf_2 _10587_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .X(_04488_));
 sky130_fd_sc_hd__inv_2 _10588_ (.A(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_1 _10589_ (.A(_04489_),
    .B(_04449_),
    .Y(_04490_));
 sky130_fd_sc_hd__inv_2 _10590_ (.A(\core.cpu_state[3] ),
    .Y(_04491_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10591_ (.A(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_2 _10592_ (.A(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__nor2_1 _10593_ (.A(_04493_),
    .B(_04378_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor3_1 _10594_ (.A(_04468_),
    .B(\core.is_sll_srl_sra ),
    .C(_04478_),
    .Y(_04495_));
 sky130_fd_sc_hd__inv_2 _10595_ (.A(_04473_),
    .Y(_04496_));
 sky130_fd_sc_hd__clkbuf_2 _10596_ (.A(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__buf_2 _10597_ (.A(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__a31o_1 _10598_ (.A1(_04472_),
    .A2(_04464_),
    .A3(_04495_),
    .B1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__a22o_1 _10599_ (.A1(_04490_),
    .A2(_04494_),
    .B1(_04499_),
    .B2(_04450_),
    .X(_00013_));
 sky130_fd_sc_hd__inv_2 _10600_ (.A(_04391_),
    .Y(_04500_));
 sky130_fd_sc_hd__inv_2 _10601_ (.A(\core.decoder_trigger ),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_2 _10602_ (.A(\core.instr_jal ),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__inv_2 _10603_ (.A(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__or3_4 _10604_ (.A(_04500_),
    .B(_04503_),
    .C(_04449_),
    .X(_04504_));
 sky130_fd_sc_hd__inv_2 _10605_ (.A(_04504_),
    .Y(_00012_));
 sky130_fd_sc_hd__nor2_2 _10606_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .B(_04492_),
    .Y(_04505_));
 sky130_fd_sc_hd__inv_2 _10607_ (.A(\core.cpu_state[4] ),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_1 _10608_ (.A(_04506_),
    .B(_04483_),
    .Y(_04507_));
 sky130_fd_sc_hd__a211o_1 _10609_ (.A1(_04391_),
    .A2(_04503_),
    .B1(_04505_),
    .C1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__nor2_1 _10610_ (.A(_04395_),
    .B(_04461_),
    .Y(_00509_));
 sky130_fd_sc_hd__a211o_1 _10611_ (.A1(_04466_),
    .A2(_04478_),
    .B1(_04508_),
    .C1(_00509_),
    .X(_04509_));
 sky130_fd_sc_hd__buf_1 _10612_ (.A(\core.cpu_state[3] ),
    .X(_04510_));
 sky130_fd_sc_hd__buf_2 _10613_ (.A(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__inv_2 _10614_ (.A(net34),
    .Y(_04512_));
 sky130_fd_sc_hd__clkbuf_2 _10615_ (.A(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_4 _10616_ (.A(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__a31o_1 _10617_ (.A1(_04490_),
    .A2(_04511_),
    .A3(_04377_),
    .B1(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__a21o_1 _10618_ (.A1(_04509_),
    .A2(_04460_),
    .B1(_04515_),
    .X(_00011_));
 sky130_fd_sc_hd__clkbuf_2 _10619_ (.A(_04440_),
    .X(_04516_));
 sky130_fd_sc_hd__or3_1 _10620_ (.A(_04384_),
    .B(_04382_),
    .C(_04381_),
    .X(_04517_));
 sky130_fd_sc_hd__a21bo_1 _10621_ (.A1(_04455_),
    .A2(_04404_),
    .B1_N(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__a21o_1 _10622_ (.A1(_04409_),
    .A2(_04516_),
    .B1(_04518_),
    .X(_00019_));
 sky130_fd_sc_hd__buf_2 _10623_ (.A(_04485_),
    .X(_04519_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10624_ (.A(_00000_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_2 _10625_ (.A(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_2 _10626_ (.A(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(\core.cpuregs[0][2] ),
    .A1(\core.cpuregs[1][2] ),
    .S(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__buf_2 _10628_ (.A(_00000_),
    .X(_04524_));
 sky130_fd_sc_hd__buf_2 _10629_ (.A(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__buf_2 _10630_ (.A(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(\core.cpuregs[2][2] ),
    .A1(\core.cpuregs[3][2] ),
    .S(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_2 _10632_ (.A(_00001_),
    .X(_04528_));
 sky130_fd_sc_hd__buf_2 _10633_ (.A(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(_04523_),
    .A1(_04527_),
    .S(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__buf_2 _10635_ (.A(_04524_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_2 _10636_ (.A(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(\core.cpuregs[6][2] ),
    .A1(\core.cpuregs[7][2] ),
    .S(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__clkbuf_4 _10638_ (.A(_04525_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(\core.cpuregs[4][2] ),
    .A1(\core.cpuregs[5][2] ),
    .S(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__inv_2 _10640_ (.A(_00001_),
    .Y(_04536_));
 sky130_fd_sc_hd__clkbuf_2 _10641_ (.A(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__mux2_1 _10642_ (.A0(_04533_),
    .A1(_04535_),
    .S(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__clkbuf_2 _10643_ (.A(_00002_),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(_04530_),
    .A1(_04538_),
    .S(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\core.cpuregs[12][2] ),
    .A1(\core.cpuregs[13][2] ),
    .S(_04532_),
    .X(_04541_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(\core.cpuregs[14][2] ),
    .A1(\core.cpuregs[15][2] ),
    .S(_04534_),
    .X(_04542_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(_04541_),
    .A1(_04542_),
    .S(_04529_),
    .X(_04543_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(\core.cpuregs[8][2] ),
    .A1(\core.cpuregs[9][2] ),
    .S(_04526_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_4 _10649_ (.A(_04525_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\core.cpuregs[10][2] ),
    .A1(\core.cpuregs[11][2] ),
    .S(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_2 _10651_ (.A(_04528_),
    .X(_04547_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(_04544_),
    .A1(_04546_),
    .S(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__inv_4 _10653_ (.A(_00002_),
    .Y(_04549_));
 sky130_fd_sc_hd__clkbuf_4 _10654_ (.A(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(_04543_),
    .A1(_04548_),
    .S(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__clkbuf_2 _10656_ (.A(_00003_),
    .X(_04552_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(_04540_),
    .A1(_04551_),
    .S(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(\core.cpuregs[16][2] ),
    .A1(\core.cpuregs[17][2] ),
    .S(_04526_),
    .X(_04554_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\core.cpuregs[18][2] ),
    .A1(\core.cpuregs[19][2] ),
    .S(_04545_),
    .X(_04555_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(_04554_),
    .A1(_04555_),
    .S(_04529_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(\core.cpuregs[22][2] ),
    .A1(\core.cpuregs[23][2] ),
    .S(_04545_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_2 _10662_ (.A(_04525_),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(\core.cpuregs[20][2] ),
    .A1(\core.cpuregs[21][2] ),
    .S(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_2 _10664_ (.A(_04536_),
    .X(_04560_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(_04557_),
    .A1(_04559_),
    .S(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(_04556_),
    .A1(_04561_),
    .S(_04539_),
    .X(_04562_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(\core.cpuregs[24][2] ),
    .A1(\core.cpuregs[25][2] ),
    .S(_04534_),
    .X(_04563_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\core.cpuregs[26][2] ),
    .A1(\core.cpuregs[27][2] ),
    .S(_04558_),
    .X(_04564_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(_04563_),
    .A1(_04564_),
    .S(_04547_),
    .X(_04565_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\core.cpuregs[28][2] ),
    .A1(\core.cpuregs[29][2] ),
    .S(_04558_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_2 _10671_ (.A(_04531_),
    .X(_04567_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\core.cpuregs[30][2] ),
    .A1(\core.cpuregs[31][2] ),
    .S(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(_04566_),
    .A1(_04568_),
    .S(_04547_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_4 _10674_ (.A(_00002_),
    .X(_04570_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(_04565_),
    .A1(_04569_),
    .S(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(_04562_),
    .A1(_04571_),
    .S(_04552_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_4 _10677_ (.A(_00004_),
    .X(_04573_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(_04553_),
    .A1(_04572_),
    .S(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10679_ (.A(\core.decoded_imm_j[3] ),
    .X(_04575_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10680_ (.A(\core.decoded_imm_j[4] ),
    .X(_04576_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10681_ (.A(\core.decoded_imm_j[11] ),
    .X(_04577_));
 sky130_fd_sc_hd__inv_2 _10682_ (.A(\core.decoded_imm_j[1] ),
    .Y(_04578_));
 sky130_fd_sc_hd__inv_2 _10683_ (.A(\core.decoded_imm_j[2] ),
    .Y(_04579_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_04578_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__or4_1 _10685_ (.A(_04575_),
    .B(_04576_),
    .C(_04577_),
    .D(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_2 _10686_ (.A(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(_04574_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _10688_ (.A(\core.decoded_imm_j[2] ),
    .B(_04519_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_1 _10689_ (.A1(_04519_),
    .A2(_04583_),
    .B1(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10690_ (.A(_04506_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_2 _10691_ (.A(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__buf_2 _10692_ (.A(_04586_),
    .X(_04588_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10693_ (.A(_04481_),
    .X(_04589_));
 sky130_fd_sc_hd__inv_2 _10694_ (.A(_04507_),
    .Y(_04590_));
 sky130_fd_sc_hd__o31a_1 _10695_ (.A1(_04588_),
    .A2(\core.reg_sh[2] ),
    .A3(_04589_),
    .B1(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__a21bo_1 _10696_ (.A1(_04585_),
    .A2(_04587_),
    .B1_N(_04591_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\core.cpuregs[0][3] ),
    .A1(\core.cpuregs[1][3] ),
    .S(_04522_),
    .X(_04592_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\core.cpuregs[2][3] ),
    .A1(\core.cpuregs[3][3] ),
    .S(_04526_),
    .X(_04593_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(_04592_),
    .A1(_04593_),
    .S(_04529_),
    .X(_04594_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\core.cpuregs[6][3] ),
    .A1(\core.cpuregs[7][3] ),
    .S(_04532_),
    .X(_04595_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\core.cpuregs[4][3] ),
    .A1(\core.cpuregs[5][3] ),
    .S(_04534_),
    .X(_04596_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(_04595_),
    .A1(_04596_),
    .S(_04560_),
    .X(_04597_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(_04594_),
    .A1(_04597_),
    .S(_04539_),
    .X(_04598_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(\core.cpuregs[12][3] ),
    .A1(\core.cpuregs[13][3] ),
    .S(_04532_),
    .X(_04599_));
 sky130_fd_sc_hd__mux2_2 _10705_ (.A0(\core.cpuregs[14][3] ),
    .A1(\core.cpuregs[15][3] ),
    .S(_04534_),
    .X(_04600_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(_04599_),
    .A1(_04600_),
    .S(_04529_),
    .X(_04601_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(\core.cpuregs[8][3] ),
    .A1(\core.cpuregs[9][3] ),
    .S(_04526_),
    .X(_04602_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\core.cpuregs[10][3] ),
    .A1(\core.cpuregs[11][3] ),
    .S(_04545_),
    .X(_04603_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(_04602_),
    .A1(_04603_),
    .S(_04547_),
    .X(_04604_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(_04601_),
    .A1(_04604_),
    .S(_04550_),
    .X(_04605_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(_04598_),
    .A1(_04605_),
    .S(_04552_),
    .X(_04606_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\core.cpuregs[16][3] ),
    .A1(\core.cpuregs[17][3] ),
    .S(_04526_),
    .X(_04607_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(\core.cpuregs[18][3] ),
    .A1(\core.cpuregs[19][3] ),
    .S(_04545_),
    .X(_04608_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(_04607_),
    .A1(_04608_),
    .S(_04529_),
    .X(_04609_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\core.cpuregs[22][3] ),
    .A1(\core.cpuregs[23][3] ),
    .S(_04545_),
    .X(_04610_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\core.cpuregs[20][3] ),
    .A1(\core.cpuregs[21][3] ),
    .S(_04558_),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(_04610_),
    .A1(_04611_),
    .S(_04560_),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(_04609_),
    .A1(_04612_),
    .S(_04539_),
    .X(_04613_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(\core.cpuregs[24][3] ),
    .A1(\core.cpuregs[25][3] ),
    .S(_04534_),
    .X(_04614_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\core.cpuregs[26][3] ),
    .A1(\core.cpuregs[27][3] ),
    .S(_04558_),
    .X(_04615_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(_04614_),
    .A1(_04615_),
    .S(_04547_),
    .X(_04616_));
 sky130_fd_sc_hd__mux2_2 _10722_ (.A0(\core.cpuregs[28][3] ),
    .A1(\core.cpuregs[29][3] ),
    .S(_04558_),
    .X(_04617_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(\core.cpuregs[30][3] ),
    .A1(\core.cpuregs[31][3] ),
    .S(_04567_),
    .X(_04618_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(_04617_),
    .A1(_04618_),
    .S(_04547_),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(_04616_),
    .A1(_04619_),
    .S(_04570_),
    .X(_04620_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(_04613_),
    .A1(_04620_),
    .S(_04552_),
    .X(_04621_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(_04606_),
    .A1(_04621_),
    .S(_04573_),
    .X(_04622_));
 sky130_fd_sc_hd__nand2_1 _10728_ (.A(_04622_),
    .B(_04582_),
    .Y(_04623_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(_04575_),
    .B(_04519_),
    .Y(_04624_));
 sky130_fd_sc_hd__o21ai_1 _10730_ (.A1(_04519_),
    .A2(_04623_),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__buf_2 _10731_ (.A(_04481_),
    .X(_04626_));
 sky130_fd_sc_hd__nor2_1 _10732_ (.A(_04506_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__nand2_1 _10733_ (.A(\core.reg_sh[3] ),
    .B(\core.reg_sh[2] ),
    .Y(_04628_));
 sky130_fd_sc_hd__nand2_1 _10734_ (.A(_04480_),
    .B(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a21o_1 _10735_ (.A1(_04627_),
    .A2(_04629_),
    .B1(_04507_),
    .X(_04630_));
 sky130_fd_sc_hd__a21o_1 _10736_ (.A1(_04625_),
    .A2(_04587_),
    .B1(_04630_),
    .X(_00035_));
 sky130_fd_sc_hd__and2_1 _10737_ (.A(_04480_),
    .B(\core.reg_sh[4] ),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_2 _10738_ (.A(\core.cpu_state[4] ),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_2 _10739_ (.A(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__buf_1 _10740_ (.A(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__a21oi_1 _10741_ (.A1(_04576_),
    .A2(_04519_),
    .B1(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__clkbuf_2 _10742_ (.A(_04531_),
    .X(_04636_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\core.cpuregs[0][4] ),
    .A1(\core.cpuregs[1][4] ),
    .S(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_2 _10744_ (.A(_04525_),
    .X(_04638_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\core.cpuregs[2][4] ),
    .A1(\core.cpuregs[3][4] ),
    .S(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_2 _10746_ (.A(_00001_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_2 _10747_ (.A(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(_04637_),
    .A1(_04639_),
    .S(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\core.cpuregs[6][4] ),
    .A1(\core.cpuregs[7][4] ),
    .S(_04636_),
    .X(_04643_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\core.cpuregs[4][4] ),
    .A1(\core.cpuregs[5][4] ),
    .S(_04638_),
    .X(_04644_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(_04643_),
    .A1(_04644_),
    .S(_04560_),
    .X(_04645_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(_04642_),
    .A1(_04645_),
    .S(_04570_),
    .X(_04646_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(\core.cpuregs[12][4] ),
    .A1(\core.cpuregs[13][4] ),
    .S(_04636_),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\core.cpuregs[14][4] ),
    .A1(\core.cpuregs[15][4] ),
    .S(_04638_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_2 _10755_ (.A(_04528_),
    .X(_04649_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(_04647_),
    .A1(_04648_),
    .S(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(\core.cpuregs[8][4] ),
    .A1(\core.cpuregs[9][4] ),
    .S(_04638_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_4 _10758_ (.A(_04525_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_1 _10759_ (.A0(\core.cpuregs[10][4] ),
    .A1(\core.cpuregs[11][4] ),
    .S(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(_04651_),
    .A1(_04653_),
    .S(_04649_),
    .X(_04654_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(_04650_),
    .A1(_04654_),
    .S(_04550_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_2 _10762_ (.A(_00003_),
    .X(_04656_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(_04646_),
    .A1(_04655_),
    .S(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\core.cpuregs[16][4] ),
    .A1(\core.cpuregs[17][4] ),
    .S(_04638_),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_2 _10765_ (.A0(\core.cpuregs[18][4] ),
    .A1(\core.cpuregs[19][4] ),
    .S(_04652_),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(_04658_),
    .A1(_04659_),
    .S(_04649_),
    .X(_04660_));
 sky130_fd_sc_hd__mux2_1 _10767_ (.A0(\core.cpuregs[22][4] ),
    .A1(\core.cpuregs[23][4] ),
    .S(_04652_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_2 _10768_ (.A(_04531_),
    .X(_04662_));
 sky130_fd_sc_hd__mux2_1 _10769_ (.A0(\core.cpuregs[20][4] ),
    .A1(\core.cpuregs[21][4] ),
    .S(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(_04661_),
    .A1(_04663_),
    .S(_04560_),
    .X(_04664_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(_04660_),
    .A1(_04664_),
    .S(_04570_),
    .X(_04665_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\core.cpuregs[24][4] ),
    .A1(\core.cpuregs[25][4] ),
    .S(_04652_),
    .X(_04666_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\core.cpuregs[26][4] ),
    .A1(\core.cpuregs[27][4] ),
    .S(_04652_),
    .X(_04667_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(_04666_),
    .A1(_04667_),
    .S(_04649_),
    .X(_04668_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\core.cpuregs[28][4] ),
    .A1(\core.cpuregs[29][4] ),
    .S(_04652_),
    .X(_04669_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(\core.cpuregs[30][4] ),
    .A1(\core.cpuregs[31][4] ),
    .S(_04662_),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(_04669_),
    .A1(_04670_),
    .S(_04649_),
    .X(_04671_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(_04668_),
    .A1(_04671_),
    .S(_04570_),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(_04665_),
    .A1(_04672_),
    .S(_04656_),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(_04657_),
    .A1(_04673_),
    .S(_04573_),
    .X(_04674_));
 sky130_fd_sc_hd__nand2_1 _10781_ (.A(_04674_),
    .B(_04582_),
    .Y(_04675_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(_04485_),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__a2bb2oi_1 _10783_ (.A1_N(_04484_),
    .A2_N(_04631_),
    .B1(_04635_),
    .B2(_04676_),
    .Y(_00036_));
 sky130_fd_sc_hd__clkbuf_2 _10784_ (.A(\core.pcpi_rs1[3] ),
    .X(_04677_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(\core.mem_la_wdata[3] ),
    .B(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_2 _10786_ (.A(\core.mem_la_wdata[3] ),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _10787_ (.A(_04679_),
    .B(_04677_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand2_4 _10788_ (.A(_04678_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__inv_2 _10789_ (.A(\core.mem_la_wdata[2] ),
    .Y(_04682_));
 sky130_fd_sc_hd__inv_2 _10790_ (.A(\core.pcpi_rs1[2] ),
    .Y(_04683_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(_04682_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _10792_ (.A(\core.mem_la_wdata[2] ),
    .B(\core.pcpi_rs1[2] ),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2_2 _10793_ (.A(_04684_),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_04681_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__inv_2 _10795_ (.A(\core.pcpi_rs1[1] ),
    .Y(_04688_));
 sky130_fd_sc_hd__inv_2 _10796_ (.A(\core.mem_la_wdata[1] ),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_1 _10797_ (.A(_04688_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_2 _10798_ (.A(\core.pcpi_rs1[1] ),
    .B(\core.mem_la_wdata[1] ),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_4 _10799_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__inv_2 _10800_ (.A(\core.pcpi_rs1[0] ),
    .Y(_04693_));
 sky130_fd_sc_hd__clkbuf_4 _10801_ (.A(\core.mem_la_wdata[0] ),
    .X(_04694_));
 sky130_fd_sc_hd__nand2_2 _10802_ (.A(_04693_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__clkbuf_2 _10803_ (.A(\core.mem_la_wdata[1] ),
    .X(_04696_));
 sky130_fd_sc_hd__nor2_1 _10804_ (.A(_04696_),
    .B(_04688_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21oi_4 _10805_ (.A1(_04692_),
    .A2(_04695_),
    .B1(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__buf_2 _10806_ (.A(\core.pcpi_rs1[2] ),
    .X(_04699_));
 sky130_fd_sc_hd__inv_2 _10807_ (.A(_04677_),
    .Y(_04700_));
 sky130_fd_sc_hd__nor2_1 _10808_ (.A(_04679_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__a31oi_2 _10809_ (.A1(_04681_),
    .A2(_04682_),
    .A3(_04699_),
    .B1(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__o21ai_4 _10810_ (.A1(_04687_),
    .A2(_04698_),
    .B1(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__or2_2 _10811_ (.A(\core.mem_la_wdata[7] ),
    .B(\core.pcpi_rs1[7] ),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_2 _10812_ (.A(\core.mem_la_wdata[7] ),
    .X(_04705_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(_04705_),
    .B(\core.pcpi_rs1[7] ),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_04704_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_2 _10815_ (.A(\core.mem_la_wdata[6] ),
    .B(\core.pcpi_rs1[6] ),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_2 _10816_ (.A(\core.mem_la_wdata[6] ),
    .X(_04709_));
 sky130_fd_sc_hd__nand2_4 _10817_ (.A(_04709_),
    .B(\core.pcpi_rs1[6] ),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_4 _10818_ (.A(_04708_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(_04707_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__inv_2 _10820_ (.A(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__buf_4 _10821_ (.A(\core.mem_la_wdata[5] ),
    .X(_04714_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_04714_),
    .B(\core.pcpi_rs1[5] ),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _10823_ (.A(\core.mem_la_wdata[5] ),
    .B(\core.pcpi_rs1[5] ),
    .Y(_04716_));
 sky130_fd_sc_hd__inv_2 _10824_ (.A(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor2_1 _10825_ (.A(_04715_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__inv_2 _10826_ (.A(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _10827_ (.A(\core.mem_la_wdata[4] ),
    .B(\core.pcpi_rs1[4] ),
    .Y(_04720_));
 sky130_fd_sc_hd__inv_2 _10828_ (.A(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__clkbuf_2 _10829_ (.A(\core.mem_la_wdata[4] ),
    .X(_04722_));
 sky130_fd_sc_hd__clkbuf_4 _10830_ (.A(\core.pcpi_rs1[4] ),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_2 _10831_ (.A(_04722_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_4 _10832_ (.A(_04721_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__and3_1 _10833_ (.A(_04713_),
    .B(_04719_),
    .C(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__nand2_2 _10834_ (.A(_04703_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__clkbuf_2 _10835_ (.A(\core.pcpi_rs1[5] ),
    .X(_04728_));
 sky130_fd_sc_hd__inv_2 _10836_ (.A(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__inv_2 _10837_ (.A(_04723_),
    .Y(_04730_));
 sky130_fd_sc_hd__nor2_1 _10838_ (.A(_04722_),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__nand2_1 _10839_ (.A(_04719_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__o21ai_2 _10840_ (.A1(_04714_),
    .A2(_04729_),
    .B1(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__clkbuf_2 _10841_ (.A(\core.pcpi_rs1[7] ),
    .X(_04734_));
 sky130_fd_sc_hd__inv_2 _10842_ (.A(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__buf_2 _10843_ (.A(_04707_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_4 _10844_ (.A(\core.pcpi_rs1[6] ),
    .X(_04737_));
 sky130_fd_sc_hd__inv_2 _10845_ (.A(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__nor2_1 _10846_ (.A(_04709_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nand2_1 _10847_ (.A(_04736_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__o21ai_1 _10848_ (.A1(_04705_),
    .A2(_04735_),
    .B1(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__a21oi_1 _10849_ (.A1(_04733_),
    .A2(_04713_),
    .B1(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_2 _10850_ (.A(_04727_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__nor2_1 _10851_ (.A(\core.pcpi_rs2[11] ),
    .B(\core.pcpi_rs1[11] ),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_1 _10852_ (.A(\core.pcpi_rs2[11] ),
    .B(\core.pcpi_rs1[11] ),
    .Y(_04745_));
 sky130_fd_sc_hd__inv_2 _10853_ (.A(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__or2_2 _10854_ (.A(_04744_),
    .B(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__or2_1 _10855_ (.A(\core.pcpi_rs2[10] ),
    .B(\core.pcpi_rs1[10] ),
    .X(_04748_));
 sky130_fd_sc_hd__nand2_2 _10856_ (.A(\core.pcpi_rs2[10] ),
    .B(\core.pcpi_rs1[10] ),
    .Y(_04749_));
 sky130_fd_sc_hd__nand2_1 _10857_ (.A(_04748_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_2 _10858_ (.A(_04747_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__clkbuf_2 _10859_ (.A(\core.pcpi_rs1[9] ),
    .X(_04752_));
 sky130_fd_sc_hd__nor2_2 _10860_ (.A(\core.pcpi_rs2[9] ),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _10861_ (.A(\core.pcpi_rs2[9] ),
    .B(\core.pcpi_rs1[9] ),
    .Y(_04754_));
 sky130_fd_sc_hd__inv_2 _10862_ (.A(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__or2_1 _10863_ (.A(_04753_),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__buf_2 _10864_ (.A(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__nor2_1 _10865_ (.A(\core.pcpi_rs2[8] ),
    .B(\core.pcpi_rs1[8] ),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _10866_ (.A(\core.pcpi_rs2[8] ),
    .B(\core.pcpi_rs1[8] ),
    .Y(_04759_));
 sky130_fd_sc_hd__inv_2 _10867_ (.A(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__or2_1 _10868_ (.A(_04758_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__nand2_1 _10869_ (.A(_04757_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _10870_ (.A(_04751_),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__or2_1 _10871_ (.A(\core.pcpi_rs2[15] ),
    .B(\core.pcpi_rs1[15] ),
    .X(_04764_));
 sky130_fd_sc_hd__nand2_2 _10872_ (.A(\core.pcpi_rs2[15] ),
    .B(\core.pcpi_rs1[15] ),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _10873_ (.A(_04764_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__or2_2 _10874_ (.A(\core.pcpi_rs2[14] ),
    .B(\core.pcpi_rs1[14] ),
    .X(_04767_));
 sky130_fd_sc_hd__nand2_4 _10875_ (.A(\core.pcpi_rs2[14] ),
    .B(\core.pcpi_rs1[14] ),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2_4 _10876_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _10877_ (.A(_04766_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__nor2_1 _10878_ (.A(\core.pcpi_rs2[13] ),
    .B(\core.pcpi_rs1[13] ),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_2 _10879_ (.A(\core.pcpi_rs2[13] ),
    .B(\core.pcpi_rs1[13] ),
    .Y(_04772_));
 sky130_fd_sc_hd__inv_2 _10880_ (.A(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__or2_1 _10881_ (.A(_04771_),
    .B(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10882_ (.A(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__or2_1 _10883_ (.A(\core.pcpi_rs2[12] ),
    .B(\core.pcpi_rs1[12] ),
    .X(_04776_));
 sky130_fd_sc_hd__nand2_2 _10884_ (.A(\core.pcpi_rs2[12] ),
    .B(\core.pcpi_rs1[12] ),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_2 _10885_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_2 _10886_ (.A(_04775_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__nor2_1 _10887_ (.A(_04770_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__and2_1 _10888_ (.A(_04763_),
    .B(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__nand2_1 _10889_ (.A(_04743_),
    .B(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__inv_2 _10890_ (.A(\core.pcpi_rs1[8] ),
    .Y(_04783_));
 sky130_fd_sc_hd__nor2_1 _10891_ (.A(\core.pcpi_rs2[8] ),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__nand2_1 _10892_ (.A(_04757_),
    .B(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__inv_2 _10893_ (.A(_04752_),
    .Y(_04786_));
 sky130_fd_sc_hd__or2_1 _10894_ (.A(\core.pcpi_rs2[9] ),
    .B(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__a21o_1 _10895_ (.A1(_04785_),
    .A2(_04787_),
    .B1(_04751_),
    .X(_04788_));
 sky130_fd_sc_hd__clkbuf_2 _10896_ (.A(_04747_),
    .X(_04789_));
 sky130_fd_sc_hd__inv_2 _10897_ (.A(\core.pcpi_rs1[10] ),
    .Y(_04790_));
 sky130_fd_sc_hd__nor2_1 _10898_ (.A(\core.pcpi_rs2[10] ),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__inv_2 _10899_ (.A(\core.pcpi_rs1[11] ),
    .Y(_04792_));
 sky130_fd_sc_hd__nor2_1 _10900_ (.A(\core.pcpi_rs2[11] ),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21oi_1 _10901_ (.A1(_04789_),
    .A2(_04791_),
    .B1(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _10902_ (.A(_04788_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__inv_2 _10903_ (.A(\core.pcpi_rs1[12] ),
    .Y(_04796_));
 sky130_fd_sc_hd__nor2_1 _10904_ (.A(\core.pcpi_rs2[12] ),
    .B(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(_04775_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__inv_2 _10906_ (.A(\core.pcpi_rs1[13] ),
    .Y(_04799_));
 sky130_fd_sc_hd__or2_1 _10907_ (.A(\core.pcpi_rs2[13] ),
    .B(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_04798_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__inv_2 _10909_ (.A(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10910_ (.A(_04766_),
    .X(_04803_));
 sky130_fd_sc_hd__inv_2 _10911_ (.A(\core.pcpi_rs1[14] ),
    .Y(_04804_));
 sky130_fd_sc_hd__nor2_1 _10912_ (.A(\core.pcpi_rs2[14] ),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__inv_2 _10913_ (.A(\core.pcpi_rs1[15] ),
    .Y(_04806_));
 sky130_fd_sc_hd__nor2_1 _10914_ (.A(\core.pcpi_rs2[15] ),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21oi_1 _10915_ (.A1(_04803_),
    .A2(_04805_),
    .B1(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__o21ai_1 _10916_ (.A1(_04770_),
    .A2(_04802_),
    .B1(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__a21oi_1 _10917_ (.A1(_04795_),
    .A2(_04780_),
    .B1(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_1 _10918_ (.A(_04782_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__buf_2 _10919_ (.A(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__inv_2 _10920_ (.A(\core.pcpi_rs2[27] ),
    .Y(_04813_));
 sky130_fd_sc_hd__inv_2 _10921_ (.A(\core.pcpi_rs1[27] ),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_1 _10922_ (.A(_04813_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(\core.pcpi_rs2[27] ),
    .B(\core.pcpi_rs1[27] ),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_2 _10924_ (.A(_04815_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__inv_2 _10925_ (.A(\core.pcpi_rs2[26] ),
    .Y(_04818_));
 sky130_fd_sc_hd__inv_2 _10926_ (.A(\core.pcpi_rs1[26] ),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _10927_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _10928_ (.A(\core.pcpi_rs2[26] ),
    .B(\core.pcpi_rs1[26] ),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_04820_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_2 _10930_ (.A(_04817_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__nor2_2 _10931_ (.A(\core.pcpi_rs2[25] ),
    .B(\core.pcpi_rs1[25] ),
    .Y(_04824_));
 sky130_fd_sc_hd__nand2_2 _10932_ (.A(\core.pcpi_rs2[25] ),
    .B(\core.pcpi_rs1[25] ),
    .Y(_04825_));
 sky130_fd_sc_hd__inv_2 _10933_ (.A(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__or2_1 _10934_ (.A(_04824_),
    .B(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_2 _10935_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__buf_2 _10936_ (.A(\core.pcpi_rs1[24] ),
    .X(_04829_));
 sky130_fd_sc_hd__nor2_1 _10937_ (.A(\core.pcpi_rs2[24] ),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__nand2_2 _10938_ (.A(\core.pcpi_rs2[24] ),
    .B(\core.pcpi_rs1[24] ),
    .Y(_04831_));
 sky130_fd_sc_hd__inv_2 _10939_ (.A(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__nor2_2 _10940_ (.A(_04830_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__inv_2 _10941_ (.A(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _10942_ (.A(_04828_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__nor2_1 _10943_ (.A(_04823_),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__inv_2 _10944_ (.A(\core.pcpi_rs2[31] ),
    .Y(_04837_));
 sky130_fd_sc_hd__inv_2 _10945_ (.A(\core.pcpi_rs1[31] ),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_2 _10946_ (.A(_04837_),
    .B(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(\core.pcpi_rs2[31] ),
    .B(\core.pcpi_rs1[31] ),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_4 _10948_ (.A(_04839_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__inv_2 _10949_ (.A(\core.pcpi_rs2[30] ),
    .Y(_04842_));
 sky130_fd_sc_hd__inv_2 _10950_ (.A(\core.pcpi_rs1[30] ),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_2 _10951_ (.A(_04842_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__clkbuf_4 _10952_ (.A(\core.pcpi_rs1[30] ),
    .X(_04845_));
 sky130_fd_sc_hd__nand2_1 _10953_ (.A(\core.pcpi_rs2[30] ),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _10954_ (.A(_04844_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _10955_ (.A(_04841_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__clkbuf_2 _10956_ (.A(\core.pcpi_rs1[28] ),
    .X(_04849_));
 sky130_fd_sc_hd__nor2_1 _10957_ (.A(\core.pcpi_rs2[28] ),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _10958_ (.A(\core.pcpi_rs2[28] ),
    .B(\core.pcpi_rs1[28] ),
    .Y(_04851_));
 sky130_fd_sc_hd__inv_2 _10959_ (.A(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nor2_1 _10960_ (.A(_04850_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__inv_2 _10961_ (.A(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(\core.pcpi_rs2[29] ),
    .B(\core.pcpi_rs1[29] ),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_2 _10963_ (.A(\core.pcpi_rs1[29] ),
    .X(_04856_));
 sky130_fd_sc_hd__nand2_1 _10964_ (.A(\core.pcpi_rs2[29] ),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_1 _10965_ (.A(_04855_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _10966_ (.A(_04854_),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__nor2_2 _10967_ (.A(_04848_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__nand2_2 _10968_ (.A(_04836_),
    .B(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _10969_ (.A(\core.pcpi_rs2[19] ),
    .B(\core.pcpi_rs1[19] ),
    .Y(_04862_));
 sky130_fd_sc_hd__nand2_1 _10970_ (.A(\core.pcpi_rs2[19] ),
    .B(\core.pcpi_rs1[19] ),
    .Y(_04863_));
 sky130_fd_sc_hd__inv_2 _10971_ (.A(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__or2_2 _10972_ (.A(_04862_),
    .B(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__nor2_2 _10973_ (.A(\core.pcpi_rs2[17] ),
    .B(\core.pcpi_rs1[17] ),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_2 _10974_ (.A(\core.pcpi_rs2[17] ),
    .B(\core.pcpi_rs1[17] ),
    .Y(_04867_));
 sky130_fd_sc_hd__inv_2 _10975_ (.A(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _10976_ (.A(_04866_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__inv_2 _10977_ (.A(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__or2_2 _10978_ (.A(\core.pcpi_rs2[16] ),
    .B(\core.pcpi_rs1[16] ),
    .X(_04871_));
 sky130_fd_sc_hd__nand2_1 _10979_ (.A(\core.pcpi_rs2[16] ),
    .B(\core.pcpi_rs1[16] ),
    .Y(_04872_));
 sky130_fd_sc_hd__nand2_2 _10980_ (.A(_04871_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__or2_1 _10981_ (.A(\core.pcpi_rs2[18] ),
    .B(\core.pcpi_rs1[18] ),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_4 _10982_ (.A(\core.pcpi_rs2[18] ),
    .B(\core.pcpi_rs1[18] ),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_2 _10983_ (.A(_04874_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__and4_2 _10984_ (.A(_04865_),
    .B(_04870_),
    .C(_04873_),
    .D(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__or2_1 _10985_ (.A(\core.pcpi_rs2[23] ),
    .B(\core.pcpi_rs1[23] ),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_2 _10986_ (.A(\core.pcpi_rs1[23] ),
    .X(_04879_));
 sky130_fd_sc_hd__nand2_1 _10987_ (.A(\core.pcpi_rs2[23] ),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_04878_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__or2_1 _10989_ (.A(\core.pcpi_rs2[22] ),
    .B(\core.pcpi_rs1[22] ),
    .X(_04882_));
 sky130_fd_sc_hd__nand2_2 _10990_ (.A(\core.pcpi_rs2[22] ),
    .B(\core.pcpi_rs1[22] ),
    .Y(_04883_));
 sky130_fd_sc_hd__nand2_1 _10991_ (.A(_04882_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_1 _10992_ (.A(_04881_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nor2_1 _10993_ (.A(\core.pcpi_rs2[20] ),
    .B(\core.pcpi_rs1[20] ),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_2 _10994_ (.A(\core.pcpi_rs2[20] ),
    .B(\core.pcpi_rs1[20] ),
    .Y(_04887_));
 sky130_fd_sc_hd__inv_2 _10995_ (.A(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__or2_4 _10996_ (.A(_04886_),
    .B(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__nor2_2 _10997_ (.A(\core.pcpi_rs2[21] ),
    .B(\core.pcpi_rs1[21] ),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_1 _10998_ (.A(\core.pcpi_rs2[21] ),
    .B(\core.pcpi_rs1[21] ),
    .Y(_04891_));
 sky130_fd_sc_hd__inv_2 _10999_ (.A(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__or2_1 _11000_ (.A(_04890_),
    .B(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__buf_1 _11001_ (.A(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__nand2_1 _11002_ (.A(_04889_),
    .B(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_2 _11003_ (.A(_04885_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _11004_ (.A(_04877_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__nor2_1 _11005_ (.A(_04861_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_1 _11006_ (.A(_04812_),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__inv_2 _11007_ (.A(_04861_),
    .Y(_04900_));
 sky130_fd_sc_hd__inv_2 _11008_ (.A(\core.pcpi_rs1[16] ),
    .Y(_04901_));
 sky130_fd_sc_hd__nor2_1 _11009_ (.A(\core.pcpi_rs2[16] ),
    .B(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_04870_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__inv_2 _11011_ (.A(\core.pcpi_rs1[17] ),
    .Y(_04904_));
 sky130_fd_sc_hd__or2_1 _11012_ (.A(\core.pcpi_rs2[17] ),
    .B(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__nand2_1 _11013_ (.A(_04903_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11014_ (.A(_04865_),
    .X(_04907_));
 sky130_fd_sc_hd__nand3_1 _11015_ (.A(_04906_),
    .B(_04907_),
    .C(_04876_),
    .Y(_04908_));
 sky130_fd_sc_hd__inv_2 _11016_ (.A(\core.pcpi_rs1[18] ),
    .Y(_04909_));
 sky130_fd_sc_hd__nor2_1 _11017_ (.A(\core.pcpi_rs2[18] ),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__inv_2 _11018_ (.A(\core.pcpi_rs1[19] ),
    .Y(_04911_));
 sky130_fd_sc_hd__nor2_1 _11019_ (.A(\core.pcpi_rs2[19] ),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__a21oi_2 _11020_ (.A1(_04865_),
    .A2(_04910_),
    .B1(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_2 _11021_ (.A(_04908_),
    .B(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(_04914_),
    .B(_04896_),
    .Y(_04915_));
 sky130_fd_sc_hd__inv_2 _11023_ (.A(\core.pcpi_rs1[21] ),
    .Y(_04916_));
 sky130_fd_sc_hd__inv_2 _11024_ (.A(\core.pcpi_rs1[20] ),
    .Y(_04917_));
 sky130_fd_sc_hd__nor2_1 _11025_ (.A(\core.pcpi_rs2[20] ),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__nand2_1 _11026_ (.A(_04894_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__o21ai_1 _11027_ (.A1(\core.pcpi_rs2[21] ),
    .A2(_04916_),
    .B1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__inv_2 _11028_ (.A(_04885_),
    .Y(_04921_));
 sky130_fd_sc_hd__inv_2 _11029_ (.A(_04879_),
    .Y(_04922_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11030_ (.A(_04881_),
    .X(_04923_));
 sky130_fd_sc_hd__inv_2 _11031_ (.A(\core.pcpi_rs1[22] ),
    .Y(_04924_));
 sky130_fd_sc_hd__nor2_1 _11032_ (.A(\core.pcpi_rs2[22] ),
    .B(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand2_1 _11033_ (.A(_04923_),
    .B(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__o21ai_1 _11034_ (.A1(\core.pcpi_rs2[23] ),
    .A2(_04922_),
    .B1(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a21oi_1 _11035_ (.A1(_04920_),
    .A2(_04921_),
    .B1(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _11036_ (.A(_04915_),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__buf_2 _11037_ (.A(_04858_),
    .X(_04930_));
 sky130_fd_sc_hd__inv_2 _11038_ (.A(_04849_),
    .Y(_04931_));
 sky130_fd_sc_hd__nor2_1 _11039_ (.A(\core.pcpi_rs2[28] ),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__inv_2 _11040_ (.A(_04856_),
    .Y(_04933_));
 sky130_fd_sc_hd__nor2_1 _11041_ (.A(\core.pcpi_rs2[29] ),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__a21oi_1 _11042_ (.A1(_04930_),
    .A2(_04932_),
    .B1(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__nor2_1 _11043_ (.A(\core.pcpi_rs2[31] ),
    .B(_04838_),
    .Y(_04936_));
 sky130_fd_sc_hd__a31o_1 _11044_ (.A1(_04841_),
    .A2(_04842_),
    .A3(_04845_),
    .B1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__o21ba_1 _11045_ (.A1(_04848_),
    .A2(_04935_),
    .B1_N(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__inv_2 _11046_ (.A(_04829_),
    .Y(_04939_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(\core.pcpi_rs2[24] ),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_2 _11048_ (.A(_04828_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__inv_2 _11049_ (.A(\core.pcpi_rs1[25] ),
    .Y(_04942_));
 sky130_fd_sc_hd__or2_1 _11050_ (.A(\core.pcpi_rs2[25] ),
    .B(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__nand2_2 _11051_ (.A(_04941_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__inv_2 _11052_ (.A(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _11053_ (.A(_04818_),
    .B(\core.pcpi_rs1[26] ),
    .Y(_04946_));
 sky130_fd_sc_hd__inv_2 _11054_ (.A(_04817_),
    .Y(_04947_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_04813_),
    .B(\core.pcpi_rs1[27] ),
    .Y(_04948_));
 sky130_fd_sc_hd__o21a_1 _11056_ (.A1(_04946_),
    .A2(_04947_),
    .B1(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__o21ai_2 _11057_ (.A1(_04823_),
    .A2(_04945_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _11058_ (.A(_04950_),
    .B(_04860_),
    .Y(_04951_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_04938_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__a21oi_1 _11060_ (.A1(_04900_),
    .A2(_04929_),
    .B1(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand3_1 _11061_ (.A(_04899_),
    .B(_04953_),
    .C(_04841_),
    .Y(_04954_));
 sky130_fd_sc_hd__inv_2 _11062_ (.A(_04936_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _11063_ (.A(_04954_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__and2_1 _11064_ (.A(_04956_),
    .B(\core.is_slti_blt_slt ),
    .X(_04957_));
 sky130_fd_sc_hd__nand2_1 _11065_ (.A(_04899_),
    .B(_04953_),
    .Y(_04958_));
 sky130_fd_sc_hd__nor2_1 _11066_ (.A(\core.pcpi_rs1[0] ),
    .B(_04694_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand2_1 _11067_ (.A(\core.pcpi_rs1[0] ),
    .B(\core.mem_la_wdata[0] ),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _11068_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__or2_1 _11069_ (.A(_04959_),
    .B(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__and4_1 _11070_ (.A(_04962_),
    .B(_04681_),
    .C(_04686_),
    .D(_04692_),
    .X(_04963_));
 sky130_fd_sc_hd__and3_1 _11071_ (.A(_04781_),
    .B(_04963_),
    .C(_04726_),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_1 _11072_ (.A(_04964_),
    .B(_04898_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _11073_ (.A(_04965_),
    .B(\core.instr_bne ),
    .Y(_04966_));
 sky130_fd_sc_hd__a21boi_1 _11074_ (.A1(_04958_),
    .A2(\core.instr_bgeu ),
    .B1_N(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand3_1 _11075_ (.A(_04954_),
    .B(\core.instr_bge ),
    .C(_04955_),
    .Y(_04968_));
 sky130_fd_sc_hd__nand2b_1 _11076_ (.A_N(_04958_),
    .B(\core.is_sltiu_bltu_sltu ),
    .Y(_04969_));
 sky130_fd_sc_hd__nand3_1 _11077_ (.A(_04967_),
    .B(_04968_),
    .C(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nor2_1 _11078_ (.A(_04957_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__or2_1 _11079_ (.A(\core.is_slti_blt_slt ),
    .B(\core.is_sltiu_bltu_sltu ),
    .X(_04972_));
 sky130_fd_sc_hd__or3b_1 _11080_ (.A(_04972_),
    .B(_04965_),
    .C_N(_04437_),
    .X(_04973_));
 sky130_fd_sc_hd__nand2_1 _11081_ (.A(_04971_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__clkbuf_2 _11082_ (.A(_04488_),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_1 _11083_ (.A(_04974_),
    .B(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_2 _11084_ (.A(_04378_),
    .B(\core.mem_do_rinst ),
    .Y(_04977_));
 sky130_fd_sc_hd__clkbuf_2 _11085_ (.A(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__clkbuf_2 _11086_ (.A(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__nor2_1 _11087_ (.A(_04493_),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__buf_1 _11088_ (.A(_04510_),
    .X(_04981_));
 sky130_fd_sc_hd__clkbuf_2 _11089_ (.A(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_4 _11090_ (.A(_04395_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_2 _11091_ (.A(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__a21oi_1 _11092_ (.A1(_04982_),
    .A2(_04984_),
    .B1(_04979_),
    .Y(_04985_));
 sky130_fd_sc_hd__a211o_1 _11093_ (.A1(_04976_),
    .A2(_04980_),
    .B1(_00509_),
    .C1(_04985_),
    .X(_00030_));
 sky130_fd_sc_hd__buf_2 _11094_ (.A(\core.instr_rdinstrh ),
    .X(_04986_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11095_ (.A(_04432_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_2 _11096_ (.A(\core.instr_rdinstr ),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_2 _11097_ (.A(\core.instr_rdcycleh ),
    .X(_04989_));
 sky130_fd_sc_hd__a22o_1 _11098_ (.A1(\core.count_instr[0] ),
    .A2(_04988_),
    .B1(_04989_),
    .B2(\core.count_cycle[32] ),
    .X(_04990_));
 sky130_fd_sc_hd__a221o_1 _11099_ (.A1(\core.count_instr[32] ),
    .A2(_04986_),
    .B1(_04987_),
    .B2(\core.count_cycle[0] ),
    .C1(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__and3_1 _11100_ (.A(_04491_),
    .B(_04506_),
    .C(_04399_),
    .X(_04992_));
 sky130_fd_sc_hd__clkbuf_2 _11101_ (.A(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__nor2_1 _11102_ (.A(\core.mem_wordsize[1] ),
    .B(\core.mem_wordsize[2] ),
    .Y(_04994_));
 sky130_fd_sc_hd__and2_1 _11103_ (.A(_04688_),
    .B(\core.mem_wordsize[2] ),
    .X(_04995_));
 sky130_fd_sc_hd__nor2_1 _11104_ (.A(_04994_),
    .B(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_04996_),
    .B(_04444_),
    .Y(_04997_));
 sky130_fd_sc_hd__clkbuf_4 _11106_ (.A(_04442_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_2 _11107_ (.A0(net31),
    .A1(net17),
    .S(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__nand2_1 _11108_ (.A(\core.mem_wordsize[1] ),
    .B(_04441_),
    .Y(_05000_));
 sky130_fd_sc_hd__inv_2 _11109_ (.A(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__clkbuf_2 _11110_ (.A(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__a22o_1 _11111_ (.A1(_04997_),
    .A2(net1),
    .B1(_04999_),
    .B2(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__nand2_1 _11112_ (.A(_04441_),
    .B(_04998_),
    .Y(_05004_));
 sky130_fd_sc_hd__inv_2 _11113_ (.A(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21oi_1 _11114_ (.A1(_04693_),
    .A2(\core.mem_wordsize[1] ),
    .B1(\core.mem_wordsize[2] ),
    .Y(_05006_));
 sky130_fd_sc_hd__inv_2 _11115_ (.A(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__a32o_1 _11116_ (.A1(_05005_),
    .A2(_04410_),
    .A3(net17),
    .B1(_05007_),
    .B2(net8),
    .X(_05008_));
 sky130_fd_sc_hd__and2_1 _11117_ (.A(_05008_),
    .B(_04998_),
    .X(_05009_));
 sky130_fd_sc_hd__or2_1 _11118_ (.A(_05003_),
    .B(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_1 _11119_ (.A(_04441_),
    .X(_05011_));
 sky130_fd_sc_hd__a22o_1 _11120_ (.A1(_04510_),
    .A2(\core.decoded_imm[0] ),
    .B1(_04633_),
    .B2(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__a221o_1 _11121_ (.A1(_04991_),
    .A2(_04993_),
    .B1(_05010_),
    .B2(_04459_),
    .C1(_05012_),
    .X(_01543_));
 sky130_fd_sc_hd__buf_2 _11122_ (.A(\core.instr_rdinstrh ),
    .X(_05013_));
 sky130_fd_sc_hd__buf_2 _11123_ (.A(_04432_),
    .X(_05014_));
 sky130_fd_sc_hd__buf_2 _11124_ (.A(\core.instr_rdinstr ),
    .X(_05015_));
 sky130_fd_sc_hd__buf_1 _11125_ (.A(\core.instr_rdcycleh ),
    .X(_05016_));
 sky130_fd_sc_hd__a22o_1 _11126_ (.A1(\core.count_instr[1] ),
    .A2(_05015_),
    .B1(_05016_),
    .B2(\core.count_cycle[33] ),
    .X(_05017_));
 sky130_fd_sc_hd__a221o_1 _11127_ (.A1(\core.count_instr[33] ),
    .A2(_05013_),
    .B1(_05014_),
    .B2(\core.count_cycle[1] ),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__buf_1 _11128_ (.A(_04992_),
    .X(_05019_));
 sky130_fd_sc_hd__inv_2 _11129_ (.A(\core.reg_pc[1] ),
    .Y(_05020_));
 sky130_fd_sc_hd__inv_2 _11130_ (.A(\core.decoded_imm[1] ),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _11131_ (.A(_05020_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_1 _11132_ (.A(\core.reg_pc[1] ),
    .B(\core.decoded_imm[1] ),
    .Y(_05023_));
 sky130_fd_sc_hd__and3_1 _11133_ (.A(_05022_),
    .B(_04510_),
    .C(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__nand2_4 _11134_ (.A(_04632_),
    .B(_04998_),
    .Y(_05025_));
 sky130_fd_sc_hd__inv_2 _11135_ (.A(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _11136_ (.A(_04440_),
    .B(_04442_),
    .Y(_05027_));
 sky130_fd_sc_hd__inv_2 _11137_ (.A(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__clkbuf_2 _11138_ (.A(_04997_),
    .X(_05029_));
 sky130_fd_sc_hd__a22o_1 _11139_ (.A1(net9),
    .A2(_05028_),
    .B1(_05029_),
    .B2(net12),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(net32),
    .A1(net18),
    .S(_04442_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_2 _11141_ (.A(_04688_),
    .X(_05032_));
 sky130_fd_sc_hd__nor2_1 _11142_ (.A(_04441_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__mux2_1 _11143_ (.A0(_05031_),
    .A1(net9),
    .S(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__and3_1 _11144_ (.A(_05034_),
    .B(_04411_),
    .C(_04444_),
    .X(_05035_));
 sky130_fd_sc_hd__o21a_1 _11145_ (.A1(_05030_),
    .A2(_05035_),
    .B1(_04459_),
    .X(_05036_));
 sky130_fd_sc_hd__a2111o_1 _11146_ (.A1(_05018_),
    .A2(_05019_),
    .B1(_05024_),
    .C1(_05026_),
    .D1(_05036_),
    .X(_01554_));
 sky130_fd_sc_hd__clkbuf_4 _11147_ (.A(_05014_),
    .X(_05037_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(_05037_),
    .B(\core.count_cycle[2] ),
    .Y(_05038_));
 sky130_fd_sc_hd__inv_2 _11149_ (.A(\core.instr_rdcycleh ),
    .Y(_05039_));
 sky130_fd_sc_hd__inv_2 _11150_ (.A(net112),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _11151_ (.A(\core.count_instr[34] ),
    .B(_04986_),
    .Y(_05041_));
 sky130_fd_sc_hd__clkbuf_2 _11152_ (.A(\core.instr_rdinstr ),
    .X(_05042_));
 sky130_fd_sc_hd__nand2_1 _11153_ (.A(\core.count_instr[2] ),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__o211a_1 _11154_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05041_),
    .C1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_2 _11155_ (.A(_05038_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__a22o_4 _11156_ (.A1(net19),
    .A2(_05002_),
    .B1(_05007_),
    .B2(net10),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_2 _11157_ (.A(_04998_),
    .X(_05047_));
 sky130_fd_sc_hd__nand2_2 _11158_ (.A(_05046_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__clkbuf_4 _11159_ (.A(_05032_),
    .X(_05049_));
 sky130_fd_sc_hd__and4_4 _11160_ (.A(_05049_),
    .B(_04411_),
    .C(_05011_),
    .D(net2),
    .X(_05050_));
 sky130_fd_sc_hd__a21oi_1 _11161_ (.A1(_05029_),
    .A2(net23),
    .B1(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_1 _11162_ (.A(_05048_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__inv_2 _11163_ (.A(\core.reg_pc[2] ),
    .Y(_05053_));
 sky130_fd_sc_hd__inv_2 _11164_ (.A(\core.decoded_imm[2] ),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_1 _11165_ (.A(_05053_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _11166_ (.A(\core.reg_pc[2] ),
    .B(\core.decoded_imm[2] ),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _11167_ (.A(_05055_),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_1 _11168_ (.A(_05023_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__inv_2 _11169_ (.A(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11170_ (.A(_05057_),
    .B(_05023_),
    .Y(_05060_));
 sky130_fd_sc_hd__a32o_1 _11171_ (.A1(_05059_),
    .A2(_04510_),
    .A3(_05060_),
    .B1(_04633_),
    .B2(_04699_),
    .X(_05061_));
 sky130_fd_sc_hd__a221o_1 _11172_ (.A1(_04993_),
    .A2(_05045_),
    .B1(_05052_),
    .B2(_04459_),
    .C1(_05061_),
    .X(_01565_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11173_ (.A(_04632_),
    .X(_05062_));
 sky130_fd_sc_hd__buf_1 _11174_ (.A(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__a22o_1 _11175_ (.A1(net20),
    .A2(_05002_),
    .B1(_05007_),
    .B2(net11),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _11176_ (.A(_05064_),
    .B(_05047_),
    .Y(_05065_));
 sky130_fd_sc_hd__and4_4 _11177_ (.A(_05049_),
    .B(_04410_),
    .C(_05011_),
    .D(net3),
    .X(_05066_));
 sky130_fd_sc_hd__a21oi_1 _11178_ (.A1(_05029_),
    .A2(net26),
    .B1(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__clkbuf_2 _11179_ (.A(_04399_),
    .X(_05068_));
 sky130_fd_sc_hd__a21oi_1 _11180_ (.A1(_05065_),
    .A2(_05067_),
    .B1(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_1 _11181_ (.A(_05059_),
    .B(_05056_),
    .Y(_05070_));
 sky130_fd_sc_hd__nor2_1 _11182_ (.A(\core.reg_pc[3] ),
    .B(\core.decoded_imm[3] ),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _11183_ (.A(\core.reg_pc[3] ),
    .B(\core.decoded_imm[3] ),
    .Y(_05072_));
 sky130_fd_sc_hd__inv_2 _11184_ (.A(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_1 _11185_ (.A(_05071_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__o21ai_1 _11186_ (.A1(_05074_),
    .A2(_05070_),
    .B1(_04981_),
    .Y(_05075_));
 sky130_fd_sc_hd__a21oi_1 _11187_ (.A1(_05070_),
    .A2(_05074_),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a22o_1 _11188_ (.A1(\core.count_instr[3] ),
    .A2(_05015_),
    .B1(_05016_),
    .B2(\core.count_cycle[35] ),
    .X(_05077_));
 sky130_fd_sc_hd__a221o_1 _11189_ (.A1(\core.count_instr[35] ),
    .A2(_05013_),
    .B1(_05014_),
    .B2(\core.count_cycle[3] ),
    .C1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__and2_1 _11190_ (.A(_05078_),
    .B(_05019_),
    .X(_05079_));
 sky130_fd_sc_hd__a2111o_1 _11191_ (.A1(_05063_),
    .A2(_04677_),
    .B1(_05069_),
    .C1(_05076_),
    .D1(_05079_),
    .X(_01568_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11192_ (.A(_04586_),
    .X(_05080_));
 sky130_fd_sc_hd__a22o_1 _11193_ (.A1(net21),
    .A2(_05002_),
    .B1(_05007_),
    .B2(net13),
    .X(_05081_));
 sky130_fd_sc_hd__nand2_1 _11194_ (.A(_05081_),
    .B(_05047_),
    .Y(_05082_));
 sky130_fd_sc_hd__clkbuf_2 _11195_ (.A(_04410_),
    .X(_05083_));
 sky130_fd_sc_hd__and4_1 _11196_ (.A(_05049_),
    .B(_05083_),
    .C(_05011_),
    .D(net4),
    .X(_05084_));
 sky130_fd_sc_hd__a21oi_1 _11197_ (.A1(_05029_),
    .A2(net27),
    .B1(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a21o_1 _11198_ (.A1(_05082_),
    .A2(_05085_),
    .B1(_05068_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_2 _11199_ (.A(_05013_),
    .X(_05087_));
 sky130_fd_sc_hd__buf_2 _11200_ (.A(_05015_),
    .X(_05088_));
 sky130_fd_sc_hd__buf_2 _11201_ (.A(_05016_),
    .X(_05089_));
 sky130_fd_sc_hd__a22o_1 _11202_ (.A1(\core.count_instr[4] ),
    .A2(_05088_),
    .B1(_05089_),
    .B2(\core.count_cycle[36] ),
    .X(_05090_));
 sky130_fd_sc_hd__a21oi_1 _11203_ (.A1(\core.count_instr[36] ),
    .A2(_05087_),
    .B1(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11204_ (.A(_05014_),
    .X(_05092_));
 sky130_fd_sc_hd__nand2_1 _11205_ (.A(_05092_),
    .B(\core.count_cycle[4] ),
    .Y(_05093_));
 sky130_fd_sc_hd__a21bo_1 _11206_ (.A1(_05091_),
    .A2(_05093_),
    .B1_N(_05019_),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _11207_ (.A(\core.reg_pc[4] ),
    .B(\core.decoded_imm[4] ),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(\core.reg_pc[4] ),
    .B(\core.decoded_imm[4] ),
    .Y(_05096_));
 sky130_fd_sc_hd__and2b_1 _11209_ (.A_N(_05095_),
    .B(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__inv_2 _11210_ (.A(_05071_),
    .Y(_05098_));
 sky130_fd_sc_hd__a21o_1 _11211_ (.A1(_05070_),
    .A2(_05098_),
    .B1(_05073_),
    .X(_05099_));
 sky130_fd_sc_hd__nor2_1 _11212_ (.A(_05097_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _11213_ (.A(_05099_),
    .B(_05097_),
    .Y(_05101_));
 sky130_fd_sc_hd__or3b_1 _11214_ (.A(_04492_),
    .B(_05100_),
    .C_N(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__o2111ai_2 _11215_ (.A1(_05080_),
    .A2(_04730_),
    .B1(_05086_),
    .C1(_05094_),
    .D1(_05102_),
    .Y(_01569_));
 sky130_fd_sc_hd__clkbuf_2 _11216_ (.A(_05019_),
    .X(_05103_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11217_ (.A(_05013_),
    .X(_05104_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11218_ (.A(_05014_),
    .X(_05105_));
 sky130_fd_sc_hd__a22o_1 _11219_ (.A1(\core.count_instr[5] ),
    .A2(_05088_),
    .B1(_05089_),
    .B2(\core.count_cycle[37] ),
    .X(_05106_));
 sky130_fd_sc_hd__a221o_1 _11220_ (.A1(\core.count_instr[37] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[5] ),
    .C1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__nor2_1 _11221_ (.A(\core.reg_pc[5] ),
    .B(\core.decoded_imm[5] ),
    .Y(_05108_));
 sky130_fd_sc_hd__nand2_1 _11222_ (.A(\core.reg_pc[5] ),
    .B(\core.decoded_imm[5] ),
    .Y(_05109_));
 sky130_fd_sc_hd__and2b_1 _11223_ (.A_N(_05108_),
    .B(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__nand2_2 _11224_ (.A(_05101_),
    .B(_05096_),
    .Y(_05111_));
 sky130_fd_sc_hd__or2_1 _11225_ (.A(_05110_),
    .B(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__nand2_1 _11226_ (.A(_05111_),
    .B(_05110_),
    .Y(_05113_));
 sky130_fd_sc_hd__and3_1 _11227_ (.A(_05112_),
    .B(_04981_),
    .C(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_2 _11228_ (.A(_04632_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _11229_ (.A1(net22),
    .A2(_05002_),
    .B1(_05007_),
    .B2(net14),
    .X(_05116_));
 sky130_fd_sc_hd__and4_1 _11230_ (.A(_05032_),
    .B(_04410_),
    .C(_05011_),
    .D(net5),
    .X(_05117_));
 sky130_fd_sc_hd__a221o_1 _11231_ (.A1(net28),
    .A2(_04997_),
    .B1(_05116_),
    .B2(_05047_),
    .C1(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_2 _11232_ (.A(_04392_),
    .X(_05119_));
 sky130_fd_sc_hd__a22o_1 _11233_ (.A1(_05115_),
    .A2(_04728_),
    .B1(_05118_),
    .B2(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__a211o_1 _11234_ (.A1(_05103_),
    .A2(_05107_),
    .B1(_05114_),
    .C1(_05120_),
    .X(_01570_));
 sky130_fd_sc_hd__nor2_1 _11235_ (.A(\core.reg_pc[6] ),
    .B(\core.decoded_imm[6] ),
    .Y(_05121_));
 sky130_fd_sc_hd__clkbuf_4 _11236_ (.A(\core.reg_pc[6] ),
    .X(_05122_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(_05122_),
    .B(\core.decoded_imm[6] ),
    .Y(_05123_));
 sky130_fd_sc_hd__and2b_1 _11238_ (.A_N(_05121_),
    .B(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__and2_1 _11239_ (.A(_05097_),
    .B(_05110_),
    .X(_05125_));
 sky130_fd_sc_hd__o21a_1 _11240_ (.A1(_05096_),
    .A2(_05108_),
    .B1(_05109_),
    .X(_05126_));
 sky130_fd_sc_hd__inv_2 _11241_ (.A(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__a21o_1 _11242_ (.A1(_05099_),
    .A2(_05125_),
    .B1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__or2_1 _11243_ (.A(_05124_),
    .B(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__nand2_1 _11244_ (.A(_05128_),
    .B(_05124_),
    .Y(_05130_));
 sky130_fd_sc_hd__a22o_1 _11245_ (.A1(\core.count_instr[38] ),
    .A2(\core.instr_rdinstrh ),
    .B1(\core.count_instr[6] ),
    .B2(_05015_),
    .X(_05131_));
 sky130_fd_sc_hd__a221o_1 _11246_ (.A1(_04989_),
    .A2(\core.count_cycle[38] ),
    .B1(_05014_),
    .B2(\core.count_cycle[6] ),
    .C1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _11247_ (.A1(_04633_),
    .A2(_04737_),
    .B1(_05132_),
    .B2(_04992_),
    .X(_05133_));
 sky130_fd_sc_hd__a22o_1 _11248_ (.A1(net24),
    .A2(_05002_),
    .B1(_05007_),
    .B2(net15),
    .X(_05134_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(_05134_),
    .B(_05047_),
    .Y(_05135_));
 sky130_fd_sc_hd__nand2_1 _11250_ (.A(_05029_),
    .B(net29),
    .Y(_05136_));
 sky130_fd_sc_hd__inv_2 _11251_ (.A(net6),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_1 _11252_ (.A(_05049_),
    .B(_04410_),
    .Y(_05138_));
 sky130_fd_sc_hd__or3_1 _11253_ (.A(_04693_),
    .B(_05137_),
    .C(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a31oi_2 _11254_ (.A1(_05135_),
    .A2(_05136_),
    .A3(_05139_),
    .B1(_05068_),
    .Y(_05140_));
 sky130_fd_sc_hd__a311o_1 _11255_ (.A1(_04982_),
    .A2(_05129_),
    .A3(_05130_),
    .B1(_05133_),
    .C1(_05140_),
    .X(_01571_));
 sky130_fd_sc_hd__clkbuf_4 _11256_ (.A(_04993_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_2 _11257_ (.A(_05016_),
    .X(_05142_));
 sky130_fd_sc_hd__a22o_1 _11258_ (.A1(\core.count_instr[7] ),
    .A2(_05042_),
    .B1(_05142_),
    .B2(\core.count_cycle[39] ),
    .X(_05143_));
 sky130_fd_sc_hd__a221o_1 _11259_ (.A1(\core.count_instr[39] ),
    .A2(_05087_),
    .B1(_05092_),
    .B2(\core.count_cycle[7] ),
    .C1(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__nor2_1 _11260_ (.A(\core.reg_pc[7] ),
    .B(\core.decoded_imm[7] ),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _11261_ (.A(\core.reg_pc[7] ),
    .B(\core.decoded_imm[7] ),
    .Y(_05146_));
 sky130_fd_sc_hd__and2b_1 _11262_ (.A_N(_05145_),
    .B(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__nand2_1 _11263_ (.A(_05130_),
    .B(_05123_),
    .Y(_05148_));
 sky130_fd_sc_hd__or2_1 _11264_ (.A(_05147_),
    .B(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_05148_),
    .B(_05147_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_1 _11266_ (.A(_04442_),
    .B(net16),
    .Y(_05151_));
 sky130_fd_sc_hd__mux2_4 _11267_ (.A0(net7),
    .A1(net25),
    .S(_04442_),
    .X(_05152_));
 sky130_fd_sc_hd__nand2_8 _11268_ (.A(_05152_),
    .B(_05001_),
    .Y(_05153_));
 sky130_fd_sc_hd__o21ai_1 _11269_ (.A1(_05006_),
    .A2(_05151_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__a21o_1 _11270_ (.A1(net30),
    .A2(_04997_),
    .B1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11271_ (.A(_04392_),
    .X(_05156_));
 sky130_fd_sc_hd__a22o_1 _11272_ (.A1(_05062_),
    .A2(_04734_),
    .B1(_05155_),
    .B2(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__a31o_1 _11273_ (.A1(_05149_),
    .A2(_04511_),
    .A3(_05150_),
    .B1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__a21o_1 _11274_ (.A1(_05141_),
    .A2(_05144_),
    .B1(_05158_),
    .X(_01572_));
 sky130_fd_sc_hd__a22o_1 _11275_ (.A1(\core.count_instr[8] ),
    .A2(_05088_),
    .B1(_05089_),
    .B2(\core.count_cycle[40] ),
    .X(_05159_));
 sky130_fd_sc_hd__a221o_1 _11276_ (.A1(\core.count_instr[40] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[8] ),
    .C1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(\core.reg_pc[8] ),
    .B(\core.decoded_imm[8] ),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(\core.reg_pc[8] ),
    .B(\core.decoded_imm[8] ),
    .Y(_05162_));
 sky130_fd_sc_hd__inv_2 _11279_ (.A(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _11280_ (.A(_05161_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__and2_1 _11281_ (.A(_05124_),
    .B(_05147_),
    .X(_05165_));
 sky130_fd_sc_hd__o21ai_1 _11282_ (.A1(_05123_),
    .A2(_05145_),
    .B1(_05146_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21o_1 _11283_ (.A1(_05165_),
    .A2(_05127_),
    .B1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__a31o_1 _11284_ (.A1(_05099_),
    .A2(_05125_),
    .A3(_05165_),
    .B1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__or2_1 _11285_ (.A(_05164_),
    .B(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__nand2_1 _11286_ (.A(_05168_),
    .B(_05164_),
    .Y(_05170_));
 sky130_fd_sc_hd__and3_1 _11287_ (.A(_05169_),
    .B(_04981_),
    .C(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__clkbuf_2 _11288_ (.A(_04994_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_4 _11289_ (.A(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_2 _11290_ (.A(_04440_),
    .X(_05174_));
 sky130_fd_sc_hd__a22o_1 _11291_ (.A1(net31),
    .A2(_05173_),
    .B1(_04999_),
    .B2(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__or2b_1 _11292_ (.A(\core.latched_is_lh ),
    .B_N(\core.latched_is_lb ),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_2 _11293_ (.A(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__nand2_2 _11294_ (.A(_05155_),
    .B(\core.latched_is_lb ),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _11295_ (.A(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__clkbuf_2 _11296_ (.A(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__a21o_1 _11297_ (.A1(_05175_),
    .A2(_05177_),
    .B1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__a22o_1 _11298_ (.A1(_05115_),
    .A2(\core.pcpi_rs1[8] ),
    .B1(_05181_),
    .B2(_05119_),
    .X(_05182_));
 sky130_fd_sc_hd__a211o_1 _11299_ (.A1(_05103_),
    .A2(_05160_),
    .B1(_05171_),
    .C1(_05182_),
    .X(_01573_));
 sky130_fd_sc_hd__a22o_1 _11300_ (.A1(\core.count_instr[9] ),
    .A2(_05088_),
    .B1(_05089_),
    .B2(\core.count_cycle[41] ),
    .X(_05183_));
 sky130_fd_sc_hd__a221o_1 _11301_ (.A1(\core.count_instr[41] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[9] ),
    .C1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__a22o_1 _11302_ (.A1(net32),
    .A2(_05172_),
    .B1(_05031_),
    .B2(_04440_),
    .X(_05185_));
 sky130_fd_sc_hd__a21o_1 _11303_ (.A1(_05177_),
    .A2(_05185_),
    .B1(_05180_),
    .X(_05186_));
 sky130_fd_sc_hd__a22o_1 _11304_ (.A1(_05115_),
    .A2(_04752_),
    .B1(_05186_),
    .B2(_05119_),
    .X(_05187_));
 sky130_fd_sc_hd__nor2_1 _11305_ (.A(\core.reg_pc[9] ),
    .B(\core.decoded_imm[9] ),
    .Y(_05188_));
 sky130_fd_sc_hd__nand2_1 _11306_ (.A(\core.reg_pc[9] ),
    .B(\core.decoded_imm[9] ),
    .Y(_05189_));
 sky130_fd_sc_hd__inv_2 _11307_ (.A(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_1 _11308_ (.A(_05188_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(_05170_),
    .B(_05162_),
    .Y(_05192_));
 sky130_fd_sc_hd__or2_1 _11310_ (.A(_05191_),
    .B(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__buf_1 _11311_ (.A(_04510_),
    .X(_05194_));
 sky130_fd_sc_hd__nand2_1 _11312_ (.A(_05192_),
    .B(_05191_),
    .Y(_05195_));
 sky130_fd_sc_hd__and3_1 _11313_ (.A(_05193_),
    .B(_05194_),
    .C(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__a211o_1 _11314_ (.A1(_05103_),
    .A2(_05184_),
    .B1(_05187_),
    .C1(_05196_),
    .X(_01574_));
 sky130_fd_sc_hd__a22o_1 _11315_ (.A1(\core.count_instr[10] ),
    .A2(_04988_),
    .B1(_05089_),
    .B2(\core.count_cycle[42] ),
    .X(_05197_));
 sky130_fd_sc_hd__a221o_1 _11316_ (.A1(\core.count_instr[42] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[10] ),
    .C1(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_4 _11317_ (.A(_04632_),
    .X(_05199_));
 sky130_fd_sc_hd__inv_2 _11318_ (.A(_04996_),
    .Y(_05200_));
 sky130_fd_sc_hd__a22o_1 _11319_ (.A1(net19),
    .A2(_05028_),
    .B1(_05200_),
    .B2(net2),
    .X(_05201_));
 sky130_fd_sc_hd__a21o_1 _11320_ (.A1(_05177_),
    .A2(_05201_),
    .B1(_05180_),
    .X(_05202_));
 sky130_fd_sc_hd__a22o_1 _11321_ (.A1(_05199_),
    .A2(\core.pcpi_rs1[10] ),
    .B1(_05202_),
    .B2(_05119_),
    .X(_05203_));
 sky130_fd_sc_hd__nor2_1 _11322_ (.A(\core.reg_pc[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _11323_ (.A(\core.reg_pc[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_05205_));
 sky130_fd_sc_hd__and2b_1 _11324_ (.A_N(_05204_),
    .B(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__and2_1 _11325_ (.A(_05164_),
    .B(_05191_),
    .X(_05207_));
 sky130_fd_sc_hd__o21a_1 _11326_ (.A1(_05162_),
    .A2(_05188_),
    .B1(_05189_),
    .X(_05208_));
 sky130_fd_sc_hd__a21bo_1 _11327_ (.A1(_05168_),
    .A2(_05207_),
    .B1_N(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__or2_1 _11328_ (.A(_05206_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_05209_),
    .B(_05206_),
    .Y(_05211_));
 sky130_fd_sc_hd__and3_1 _11330_ (.A(_05210_),
    .B(_05194_),
    .C(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__a211o_1 _11331_ (.A1(_05103_),
    .A2(_05198_),
    .B1(_05203_),
    .C1(_05212_),
    .X(_01544_));
 sky130_fd_sc_hd__a22o_1 _11332_ (.A1(\core.count_instr[11] ),
    .A2(_05042_),
    .B1(_05142_),
    .B2(\core.count_cycle[43] ),
    .X(_05213_));
 sky130_fd_sc_hd__a221o_1 _11333_ (.A1(\core.count_instr[43] ),
    .A2(_05087_),
    .B1(_05092_),
    .B2(\core.count_cycle[11] ),
    .C1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(\core.reg_pc[11] ),
    .B(\core.decoded_imm[11] ),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_1 _11335_ (.A(\core.reg_pc[11] ),
    .B(\core.decoded_imm[11] ),
    .Y(_05216_));
 sky130_fd_sc_hd__inv_2 _11336_ (.A(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nor2_1 _11337_ (.A(_05215_),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand2_1 _11338_ (.A(_05211_),
    .B(_05205_),
    .Y(_05219_));
 sky130_fd_sc_hd__or2_1 _11339_ (.A(_05218_),
    .B(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(_05219_),
    .B(_05218_),
    .Y(_05221_));
 sky130_fd_sc_hd__a22o_1 _11341_ (.A1(net20),
    .A2(_05028_),
    .B1(_05200_),
    .B2(net3),
    .X(_05222_));
 sky130_fd_sc_hd__a21o_1 _11342_ (.A1(_05176_),
    .A2(_05222_),
    .B1(_05179_),
    .X(_05223_));
 sky130_fd_sc_hd__a22o_1 _11343_ (.A1(_05062_),
    .A2(\core.pcpi_rs1[11] ),
    .B1(_05223_),
    .B2(_05156_),
    .X(_05224_));
 sky130_fd_sc_hd__a31o_1 _11344_ (.A1(_05220_),
    .A2(_04511_),
    .A3(_05221_),
    .B1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__a21o_1 _11345_ (.A1(_05141_),
    .A2(_05214_),
    .B1(_05225_),
    .X(_01545_));
 sky130_fd_sc_hd__a22o_1 _11346_ (.A1(\core.count_instr[12] ),
    .A2(_04988_),
    .B1(_04989_),
    .B2(\core.count_cycle[44] ),
    .X(_05226_));
 sky130_fd_sc_hd__a221o_1 _11347_ (.A1(\core.count_instr[44] ),
    .A2(_04986_),
    .B1(_04987_),
    .B2(\core.count_cycle[12] ),
    .C1(_05226_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(net21),
    .A2(_05028_),
    .B1(_05200_),
    .B2(net4),
    .X(_05228_));
 sky130_fd_sc_hd__a21o_1 _11349_ (.A1(_05177_),
    .A2(_05228_),
    .B1(_05180_),
    .X(_05229_));
 sky130_fd_sc_hd__a22o_1 _11350_ (.A1(_05199_),
    .A2(\core.pcpi_rs1[12] ),
    .B1(_05229_),
    .B2(_05119_),
    .X(_05230_));
 sky130_fd_sc_hd__nor2_1 _11351_ (.A(\core.reg_pc[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _11352_ (.A(\core.reg_pc[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_05232_));
 sky130_fd_sc_hd__and2b_1 _11353_ (.A_N(_05231_),
    .B(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__nand2_4 _11354_ (.A(_05206_),
    .B(_05218_),
    .Y(_05234_));
 sky130_fd_sc_hd__inv_2 _11355_ (.A(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__o221ai_4 _11356_ (.A1(_05205_),
    .A2(_05215_),
    .B1(_05234_),
    .B2(_05208_),
    .C1(_05216_),
    .Y(_05236_));
 sky130_fd_sc_hd__a31o_1 _11357_ (.A1(_05168_),
    .A2(_05207_),
    .A3(_05235_),
    .B1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__or2_1 _11358_ (.A(_05233_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(_05237_),
    .B(_05233_),
    .Y(_05239_));
 sky130_fd_sc_hd__and3_1 _11360_ (.A(_05238_),
    .B(_05194_),
    .C(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__a211o_1 _11361_ (.A1(_05103_),
    .A2(_05227_),
    .B1(_05230_),
    .C1(_05240_),
    .X(_01546_));
 sky130_fd_sc_hd__a22o_1 _11362_ (.A1(\core.count_instr[13] ),
    .A2(_04988_),
    .B1(_04989_),
    .B2(\core.count_cycle[45] ),
    .X(_05241_));
 sky130_fd_sc_hd__a221o_2 _11363_ (.A1(\core.count_instr[45] ),
    .A2(_04986_),
    .B1(_04987_),
    .B2(\core.count_cycle[13] ),
    .C1(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__o21ai_1 _11364_ (.A1(net22),
    .A2(_05032_),
    .B1(_05174_),
    .Y(_05243_));
 sky130_fd_sc_hd__inv_2 _11365_ (.A(_05172_),
    .Y(_05244_));
 sky130_fd_sc_hd__nand2_1 _11366_ (.A(_05243_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__a21o_1 _11367_ (.A1(_05244_),
    .A2(_04998_),
    .B1(net5),
    .X(_05246_));
 sky130_fd_sc_hd__a31o_1 _11368_ (.A1(_05177_),
    .A2(_05245_),
    .A3(_05246_),
    .B1(_05180_),
    .X(_05247_));
 sky130_fd_sc_hd__a22o_1 _11369_ (.A1(_05199_),
    .A2(\core.pcpi_rs1[13] ),
    .B1(_05247_),
    .B2(_05119_),
    .X(_05248_));
 sky130_fd_sc_hd__nor2_1 _11370_ (.A(\core.reg_pc[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_05249_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(\core.reg_pc[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_05250_));
 sky130_fd_sc_hd__or2b_2 _11372_ (.A(_05249_),
    .B_N(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__nand2_2 _11373_ (.A(_05239_),
    .B(_05232_),
    .Y(_05252_));
 sky130_fd_sc_hd__xor2_4 _11374_ (.A(_05251_),
    .B(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__nor2_1 _11375_ (.A(_04493_),
    .B(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a211o_1 _11376_ (.A1(_05103_),
    .A2(_05242_),
    .B1(_05248_),
    .C1(_05254_),
    .X(_01547_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(\core.reg_pc[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_4 _11378_ (.A(\core.reg_pc[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_05256_));
 sky130_fd_sc_hd__and2b_1 _11379_ (.A_N(_05255_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__inv_2 _11380_ (.A(_05251_),
    .Y(_05258_));
 sky130_fd_sc_hd__nand2_1 _11381_ (.A(_05258_),
    .B(_05233_),
    .Y(_05259_));
 sky130_fd_sc_hd__or2b_1 _11382_ (.A(_05259_),
    .B_N(_05237_),
    .X(_05260_));
 sky130_fd_sc_hd__o21a_1 _11383_ (.A1(_05232_),
    .A2(_05249_),
    .B1(_05250_),
    .X(_05261_));
 sky130_fd_sc_hd__nand2_1 _11384_ (.A(_05260_),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__or2_2 _11385_ (.A(_05257_),
    .B(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__nand2_2 _11386_ (.A(_05262_),
    .B(_05257_),
    .Y(_05264_));
 sky130_fd_sc_hd__nand2_1 _11387_ (.A(_05263_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__a22o_1 _11388_ (.A1(\core.count_instr[14] ),
    .A2(_05088_),
    .B1(_05089_),
    .B2(\core.count_cycle[46] ),
    .X(_05266_));
 sky130_fd_sc_hd__a221o_2 _11389_ (.A1(\core.count_instr[46] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[14] ),
    .C1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__buf_4 _11390_ (.A(_05019_),
    .X(_05268_));
 sky130_fd_sc_hd__nand2_8 _11391_ (.A(_05267_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_1 _11392_ (.A1(net24),
    .A2(_05032_),
    .B1(_05174_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_1 _11393_ (.A(_05270_),
    .B(_05244_),
    .Y(_05271_));
 sky130_fd_sc_hd__o21ai_1 _11394_ (.A1(_05049_),
    .A2(_05173_),
    .B1(_05137_),
    .Y(_05272_));
 sky130_fd_sc_hd__a31o_1 _11395_ (.A1(_05177_),
    .A2(_05271_),
    .A3(_05272_),
    .B1(_05180_),
    .X(_05273_));
 sky130_fd_sc_hd__o2bb2a_1 _11396_ (.A1_N(_04459_),
    .A2_N(_05273_),
    .B1(_05080_),
    .B2(_04804_),
    .X(_05274_));
 sky130_fd_sc_hd__o211ai_2 _11397_ (.A1(_04493_),
    .A2(_05265_),
    .B1(_05269_),
    .C1(_05274_),
    .Y(_01548_));
 sky130_fd_sc_hd__clkbuf_2 _11398_ (.A(\core.reg_pc[15] ),
    .X(_05275_));
 sky130_fd_sc_hd__nor2_2 _11399_ (.A(_05275_),
    .B(\core.decoded_imm[15] ),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_2 _11400_ (.A(\core.reg_pc[15] ),
    .B(\core.decoded_imm[15] ),
    .Y(_05277_));
 sky130_fd_sc_hd__inv_2 _11401_ (.A(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__nor2_4 _11402_ (.A(_05276_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__inv_2 _11403_ (.A(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__a21oi_4 _11404_ (.A1(_05264_),
    .A2(_05256_),
    .B1(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand3_2 _11405_ (.A(_05264_),
    .B(_05256_),
    .C(_05280_),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_8 _11406_ (.A(_05282_),
    .B(_04511_),
    .Y(_05283_));
 sky130_fd_sc_hd__or2_2 _11407_ (.A(\core.latched_is_lh ),
    .B(\core.latched_is_lb ),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_2 _11408_ (.A(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_2 _11409_ (.A(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__a22o_1 _11410_ (.A1(net7),
    .A2(_04994_),
    .B1(_05152_),
    .B2(_04440_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _11411_ (.A1(_05286_),
    .A2(_05287_),
    .B1(_04459_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand2_1 _11412_ (.A(_05287_),
    .B(\core.latched_is_lh ),
    .Y(_05289_));
 sky130_fd_sc_hd__and3_1 _11413_ (.A(_05178_),
    .B(_05284_),
    .C(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__buf_2 _11414_ (.A(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_2 _11415_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__o22a_1 _11416_ (.A1(_05080_),
    .A2(_04806_),
    .B1(_05288_),
    .B2(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_4 _11417_ (.A(_05013_),
    .X(_05294_));
 sky130_fd_sc_hd__buf_2 _11418_ (.A(_05015_),
    .X(_05295_));
 sky130_fd_sc_hd__buf_2 _11419_ (.A(_05016_),
    .X(_05296_));
 sky130_fd_sc_hd__a22o_1 _11420_ (.A1(\core.count_instr[15] ),
    .A2(_05295_),
    .B1(_05296_),
    .B2(\core.count_cycle[47] ),
    .X(_05297_));
 sky130_fd_sc_hd__a221o_1 _11421_ (.A1(\core.count_instr[47] ),
    .A2(_05294_),
    .B1(_05037_),
    .B2(\core.count_cycle[15] ),
    .C1(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__nand2_1 _11422_ (.A(_05298_),
    .B(_05268_),
    .Y(_05299_));
 sky130_fd_sc_hd__o211ai_2 _11423_ (.A1(_05281_),
    .A2(_05283_),
    .B1(_05293_),
    .C1(_05299_),
    .Y(_01549_));
 sky130_fd_sc_hd__a22o_1 _11424_ (.A1(\core.count_instr[16] ),
    .A2(_05042_),
    .B1(_05142_),
    .B2(\core.count_cycle[48] ),
    .X(_05300_));
 sky130_fd_sc_hd__a221o_1 _11425_ (.A1(\core.count_instr[48] ),
    .A2(_05087_),
    .B1(_05092_),
    .B2(\core.count_cycle[16] ),
    .C1(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__nor2_1 _11426_ (.A(\core.reg_pc[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_1 _11427_ (.A(\core.reg_pc[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_05303_));
 sky130_fd_sc_hd__inv_2 _11428_ (.A(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__nor2_1 _11429_ (.A(_05302_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _11430_ (.A(_05257_),
    .B(_05279_),
    .Y(_05306_));
 sky130_fd_sc_hd__nor2_1 _11431_ (.A(_05306_),
    .B(_05259_),
    .Y(_05307_));
 sky130_fd_sc_hd__and3_1 _11432_ (.A(_05307_),
    .B(_05207_),
    .C(_05235_),
    .X(_05308_));
 sky130_fd_sc_hd__nand2_2 _11433_ (.A(_05168_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__o221a_1 _11434_ (.A1(_05256_),
    .A2(_05280_),
    .B1(_05261_),
    .B2(_05306_),
    .C1(_05277_),
    .X(_05310_));
 sky130_fd_sc_hd__a21boi_4 _11435_ (.A1(_05236_),
    .A2(_05307_),
    .B1_N(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__nand2_4 _11436_ (.A(_05309_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__nor2_1 _11437_ (.A(_05305_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_1 _11438_ (.A(_05312_),
    .B(_05305_),
    .Y(_05314_));
 sky130_fd_sc_hd__or3b_2 _11439_ (.A(_04492_),
    .B(_05313_),
    .C_N(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_2 _11440_ (.A(_04399_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_2 _11441_ (.A(_05173_),
    .X(_05317_));
 sky130_fd_sc_hd__a21oi_1 _11442_ (.A1(_05317_),
    .A2(net8),
    .B1(_05285_),
    .Y(_05318_));
 sky130_fd_sc_hd__clkbuf_2 _11443_ (.A(_04586_),
    .X(_05319_));
 sky130_fd_sc_hd__o32a_2 _11444_ (.A1(_05316_),
    .A2(_05318_),
    .A3(_05291_),
    .B1(_05319_),
    .B2(_04901_),
    .X(_05320_));
 sky130_fd_sc_hd__nand2_4 _11445_ (.A(_05315_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__a21o_1 _11446_ (.A1(_05141_),
    .A2(_05301_),
    .B1(_05321_),
    .X(_01550_));
 sky130_fd_sc_hd__a22o_1 _11447_ (.A1(\core.count_instr[17] ),
    .A2(_05042_),
    .B1(_05142_),
    .B2(\core.count_cycle[49] ),
    .X(_05322_));
 sky130_fd_sc_hd__a221o_1 _11448_ (.A1(\core.count_instr[49] ),
    .A2(_05087_),
    .B1(_05092_),
    .B2(\core.count_cycle[17] ),
    .C1(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__nor2_1 _11449_ (.A(\core.reg_pc[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_1 _11450_ (.A(\core.reg_pc[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_05325_));
 sky130_fd_sc_hd__and2b_1 _11451_ (.A_N(_05324_),
    .B(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__nand2_1 _11452_ (.A(_05314_),
    .B(_05303_),
    .Y(_05327_));
 sky130_fd_sc_hd__or2_1 _11453_ (.A(_05326_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__nand2_1 _11454_ (.A(_05327_),
    .B(_05326_),
    .Y(_05329_));
 sky130_fd_sc_hd__a21oi_1 _11455_ (.A1(_05173_),
    .A2(net9),
    .B1(_05285_),
    .Y(_05330_));
 sky130_fd_sc_hd__nor2_1 _11456_ (.A(_05330_),
    .B(_05291_),
    .Y(_05331_));
 sky130_fd_sc_hd__a22o_1 _11457_ (.A1(_05062_),
    .A2(\core.pcpi_rs1[17] ),
    .B1(_05331_),
    .B2(_05156_),
    .X(_05332_));
 sky130_fd_sc_hd__a31o_1 _11458_ (.A1(_05328_),
    .A2(_04511_),
    .A3(_05329_),
    .B1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a21o_1 _11459_ (.A1(_05141_),
    .A2(_05323_),
    .B1(_05333_),
    .X(_01551_));
 sky130_fd_sc_hd__a22o_1 _11460_ (.A1(\core.count_instr[18] ),
    .A2(_04988_),
    .B1(_04989_),
    .B2(\core.count_cycle[50] ),
    .X(_05334_));
 sky130_fd_sc_hd__a221o_1 _11461_ (.A1(\core.count_instr[50] ),
    .A2(_04986_),
    .B1(_04987_),
    .B2(\core.count_cycle[18] ),
    .C1(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__a21oi_1 _11462_ (.A1(_05317_),
    .A2(net10),
    .B1(_05285_),
    .Y(_05336_));
 sky130_fd_sc_hd__nor2_4 _11463_ (.A(_05336_),
    .B(_05291_),
    .Y(_05337_));
 sky130_fd_sc_hd__a22o_1 _11464_ (.A1(_05199_),
    .A2(\core.pcpi_rs1[18] ),
    .B1(_05337_),
    .B2(_05156_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_4 _11465_ (.A(\core.reg_pc[18] ),
    .X(_05339_));
 sky130_fd_sc_hd__nor2_1 _11466_ (.A(_05339_),
    .B(\core.decoded_imm[18] ),
    .Y(_05340_));
 sky130_fd_sc_hd__nand2_2 _11467_ (.A(_05339_),
    .B(\core.decoded_imm[18] ),
    .Y(_05341_));
 sky130_fd_sc_hd__and2b_1 _11468_ (.A_N(_05340_),
    .B(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__nand2_2 _11469_ (.A(_05326_),
    .B(_05305_),
    .Y(_05343_));
 sky130_fd_sc_hd__inv_2 _11470_ (.A(_05312_),
    .Y(_05344_));
 sky130_fd_sc_hd__o21a_1 _11471_ (.A1(_05303_),
    .A2(_05324_),
    .B1(_05325_),
    .X(_05345_));
 sky130_fd_sc_hd__o21ai_2 _11472_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(_05342_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__nand2_1 _11474_ (.A(_05346_),
    .B(_05342_),
    .Y(_05348_));
 sky130_fd_sc_hd__and3_1 _11475_ (.A(_05347_),
    .B(_05194_),
    .C(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__a211o_1 _11476_ (.A1(_04993_),
    .A2(_05335_),
    .B1(_05338_),
    .C1(_05349_),
    .X(_01552_));
 sky130_fd_sc_hd__clkbuf_2 _11477_ (.A(_05013_),
    .X(_05350_));
 sky130_fd_sc_hd__buf_2 _11478_ (.A(_05015_),
    .X(_05351_));
 sky130_fd_sc_hd__a22o_1 _11479_ (.A1(\core.count_instr[19] ),
    .A2(_05351_),
    .B1(_05142_),
    .B2(\core.count_cycle[51] ),
    .X(_05352_));
 sky130_fd_sc_hd__a221o_1 _11480_ (.A1(\core.count_instr[51] ),
    .A2(_05350_),
    .B1(_05092_),
    .B2(\core.count_cycle[19] ),
    .C1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_4 _11481_ (.A(_04493_),
    .X(_05354_));
 sky130_fd_sc_hd__nor2_1 _11482_ (.A(\core.reg_pc[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_2 _11483_ (.A(\core.reg_pc[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_05356_));
 sky130_fd_sc_hd__inv_2 _11484_ (.A(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__nor2_1 _11485_ (.A(_05355_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__inv_2 _11486_ (.A(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__nand2_1 _11487_ (.A(_05348_),
    .B(_05341_),
    .Y(_05360_));
 sky130_fd_sc_hd__xor2_1 _11488_ (.A(_05359_),
    .B(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11489_ (.A(_04399_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_2 _11490_ (.A(_05173_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_2 _11491_ (.A(_05284_),
    .X(_05364_));
 sky130_fd_sc_hd__a21oi_1 _11492_ (.A1(_05363_),
    .A2(net11),
    .B1(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__clkbuf_4 _11493_ (.A(_05290_),
    .X(_05366_));
 sky130_fd_sc_hd__o32a_1 _11494_ (.A1(_05362_),
    .A2(_05365_),
    .A3(_05366_),
    .B1(_05080_),
    .B2(_04911_),
    .X(_05367_));
 sky130_fd_sc_hd__o21ai_1 _11495_ (.A1(_05354_),
    .A2(_05361_),
    .B1(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__a21o_1 _11496_ (.A1(_05141_),
    .A2(_05353_),
    .B1(_05368_),
    .X(_01553_));
 sky130_fd_sc_hd__a22o_1 _11497_ (.A1(\core.count_instr[20] ),
    .A2(_04988_),
    .B1(_04989_),
    .B2(\core.count_cycle[52] ),
    .X(_05369_));
 sky130_fd_sc_hd__a221o_1 _11498_ (.A1(\core.count_instr[52] ),
    .A2(_04986_),
    .B1(_04987_),
    .B2(\core.count_cycle[20] ),
    .C1(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a21oi_2 _11499_ (.A1(_05317_),
    .A2(net13),
    .B1(_05285_),
    .Y(_05371_));
 sky130_fd_sc_hd__nor2_4 _11500_ (.A(_05371_),
    .B(_05291_),
    .Y(_05372_));
 sky130_fd_sc_hd__a22o_1 _11501_ (.A1(_05199_),
    .A2(\core.pcpi_rs1[20] ),
    .B1(_05372_),
    .B2(_05156_),
    .X(_05373_));
 sky130_fd_sc_hd__nor2_1 _11502_ (.A(\core.reg_pc[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_05374_));
 sky130_fd_sc_hd__nand2_2 _11503_ (.A(\core.reg_pc[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_05375_));
 sky130_fd_sc_hd__and2b_1 _11504_ (.A_N(_05374_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__nand2_1 _11505_ (.A(_05342_),
    .B(_05358_),
    .Y(_05377_));
 sky130_fd_sc_hd__nor2_1 _11506_ (.A(_05343_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__o221a_1 _11507_ (.A1(_05341_),
    .A2(_05359_),
    .B1(_05345_),
    .B2(_05377_),
    .C1(_05356_),
    .X(_05379_));
 sky130_fd_sc_hd__a21bo_1 _11508_ (.A1(_05312_),
    .A2(_05378_),
    .B1_N(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__or2_1 _11509_ (.A(_05376_),
    .B(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__nand2_1 _11510_ (.A(_05380_),
    .B(_05376_),
    .Y(_05382_));
 sky130_fd_sc_hd__and3_1 _11511_ (.A(_05381_),
    .B(_04981_),
    .C(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__a211o_1 _11512_ (.A1(_04993_),
    .A2(_05370_),
    .B1(_05373_),
    .C1(_05383_),
    .X(_01555_));
 sky130_fd_sc_hd__clkbuf_2 _11513_ (.A(_04987_),
    .X(_05384_));
 sky130_fd_sc_hd__buf_2 _11514_ (.A(_05016_),
    .X(_05385_));
 sky130_fd_sc_hd__a22o_1 _11515_ (.A1(\core.count_instr[21] ),
    .A2(_05351_),
    .B1(_05385_),
    .B2(\core.count_cycle[53] ),
    .X(_05386_));
 sky130_fd_sc_hd__a221o_1 _11516_ (.A1(\core.count_instr[53] ),
    .A2(_05350_),
    .B1(_05384_),
    .B2(\core.count_cycle[21] ),
    .C1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__nor2_1 _11517_ (.A(\core.reg_pc[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _11518_ (.A(\core.reg_pc[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_05389_));
 sky130_fd_sc_hd__and2b_1 _11519_ (.A_N(_05388_),
    .B(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_05382_),
    .B(_05375_),
    .Y(_05391_));
 sky130_fd_sc_hd__or2_1 _11521_ (.A(_05390_),
    .B(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__nand2_1 _11522_ (.A(_05391_),
    .B(_05390_),
    .Y(_05393_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_05392_),
    .B(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__a21oi_1 _11524_ (.A1(_05363_),
    .A2(net14),
    .B1(_05364_),
    .Y(_05395_));
 sky130_fd_sc_hd__o32a_1 _11525_ (.A1(_05362_),
    .A2(_05395_),
    .A3(_05366_),
    .B1(_05080_),
    .B2(_04916_),
    .X(_05396_));
 sky130_fd_sc_hd__o21ai_1 _11526_ (.A1(_05354_),
    .A2(_05394_),
    .B1(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a21o_1 _11527_ (.A1(_05141_),
    .A2(_05387_),
    .B1(_05397_),
    .X(_01556_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11528_ (.A(_05019_),
    .X(_05398_));
 sky130_fd_sc_hd__a22o_1 _11529_ (.A1(\core.count_instr[22] ),
    .A2(_05351_),
    .B1(_05385_),
    .B2(\core.count_cycle[54] ),
    .X(_05399_));
 sky130_fd_sc_hd__a221o_1 _11530_ (.A1(\core.count_instr[54] ),
    .A2(_05350_),
    .B1(_05384_),
    .B2(\core.count_cycle[22] ),
    .C1(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__nor2_1 _11531_ (.A(\core.reg_pc[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_05401_));
 sky130_fd_sc_hd__nand2_2 _11532_ (.A(\core.reg_pc[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_05402_));
 sky130_fd_sc_hd__inv_2 _11533_ (.A(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__or2_1 _11534_ (.A(_05401_),
    .B(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__inv_2 _11535_ (.A(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(_05376_),
    .B(_05390_),
    .Y(_05406_));
 sky130_fd_sc_hd__inv_2 _11537_ (.A(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _11538_ (.A(_05380_),
    .B(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__o21a_1 _11539_ (.A1(_05375_),
    .A2(_05388_),
    .B1(_05389_),
    .X(_05409_));
 sky130_fd_sc_hd__nand2_1 _11540_ (.A(_05408_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__or2_1 _11541_ (.A(_05405_),
    .B(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__nand2_1 _11542_ (.A(_05410_),
    .B(_05405_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__a21oi_2 _11544_ (.A1(_05363_),
    .A2(net15),
    .B1(_05364_),
    .Y(_05414_));
 sky130_fd_sc_hd__o32a_1 _11545_ (.A1(_05362_),
    .A2(_05414_),
    .A3(_05366_),
    .B1(_05319_),
    .B2(_04924_),
    .X(_05415_));
 sky130_fd_sc_hd__o21ai_2 _11546_ (.A1(_05354_),
    .A2(_05413_),
    .B1(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21o_1 _11547_ (.A1(_05398_),
    .A2(_05400_),
    .B1(_05416_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _11548_ (.A(\core.reg_pc[23] ),
    .B(\core.decoded_imm[23] ),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _11549_ (.A(\core.reg_pc[23] ),
    .B(\core.decoded_imm[23] ),
    .Y(_05418_));
 sky130_fd_sc_hd__and2b_1 _11550_ (.A_N(_05417_),
    .B(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(_05412_),
    .B(_05402_),
    .Y(_05420_));
 sky130_fd_sc_hd__or2_2 _11552_ (.A(_05419_),
    .B(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__nand2_1 _11553_ (.A(_05420_),
    .B(_05419_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand3_2 _11554_ (.A(_05421_),
    .B(_04982_),
    .C(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__clkbuf_2 _11555_ (.A(_05172_),
    .X(_05424_));
 sky130_fd_sc_hd__a21oi_1 _11556_ (.A1(_05424_),
    .A2(net16),
    .B1(_05286_),
    .Y(_05425_));
 sky130_fd_sc_hd__o32a_1 _11557_ (.A1(_05068_),
    .A2(_05425_),
    .A3(_05292_),
    .B1(_04587_),
    .B2(_04922_),
    .X(_05426_));
 sky130_fd_sc_hd__a22o_1 _11558_ (.A1(\core.count_instr[23] ),
    .A2(_05295_),
    .B1(_05296_),
    .B2(\core.count_cycle[55] ),
    .X(_05427_));
 sky130_fd_sc_hd__a221o_1 _11559_ (.A1(\core.count_instr[55] ),
    .A2(_05294_),
    .B1(_05037_),
    .B2(\core.count_cycle[23] ),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_05428_),
    .B(_05398_),
    .Y(_05429_));
 sky130_fd_sc_hd__nand3_1 _11561_ (.A(_05423_),
    .B(_05426_),
    .C(_05429_),
    .Y(_01558_));
 sky130_fd_sc_hd__a22o_1 _11562_ (.A1(\core.count_instr[24] ),
    .A2(_05351_),
    .B1(_05385_),
    .B2(\core.count_cycle[56] ),
    .X(_05430_));
 sky130_fd_sc_hd__a221o_1 _11563_ (.A1(\core.count_instr[56] ),
    .A2(_05350_),
    .B1(_05384_),
    .B2(\core.count_cycle[24] ),
    .C1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_1 _11564_ (.A(\core.reg_pc[24] ),
    .B(\core.decoded_imm[24] ),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_2 _11565_ (.A(\core.reg_pc[24] ),
    .B(\core.decoded_imm[24] ),
    .Y(_05433_));
 sky130_fd_sc_hd__inv_2 _11566_ (.A(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__nor2_2 _11567_ (.A(_05432_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__and2_1 _11568_ (.A(_05405_),
    .B(_05419_),
    .X(_05436_));
 sky130_fd_sc_hd__and3_1 _11569_ (.A(_05436_),
    .B(_05378_),
    .C(_05407_),
    .X(_05437_));
 sky130_fd_sc_hd__nand2_1 _11570_ (.A(_05312_),
    .B(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(_05436_),
    .B(_05407_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_05419_),
    .B(_05403_),
    .Y(_05440_));
 sky130_fd_sc_hd__o311a_1 _11573_ (.A1(_05417_),
    .A2(_05404_),
    .A3(_05409_),
    .B1(_05418_),
    .C1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__o21a_1 _11574_ (.A1(_05379_),
    .A2(_05439_),
    .B1(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__nand2_2 _11575_ (.A(_05438_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__or2_1 _11576_ (.A(_05435_),
    .B(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__nand2_1 _11577_ (.A(_05443_),
    .B(_05435_),
    .Y(_05445_));
 sky130_fd_sc_hd__a21oi_2 _11578_ (.A1(_05173_),
    .A2(net17),
    .B1(_05285_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_1 _11579_ (.A(_05446_),
    .B(_05291_),
    .Y(_05447_));
 sky130_fd_sc_hd__a22o_1 _11580_ (.A1(_05062_),
    .A2(_04829_),
    .B1(_05447_),
    .B2(_05156_),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _11581_ (.A1(_05444_),
    .A2(_05194_),
    .A3(_05445_),
    .B1(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__a21o_1 _11582_ (.A1(_05398_),
    .A2(_05431_),
    .B1(_05449_),
    .X(_01559_));
 sky130_fd_sc_hd__a22o_1 _11583_ (.A1(\core.count_instr[25] ),
    .A2(_05351_),
    .B1(_05385_),
    .B2(\core.count_cycle[57] ),
    .X(_05450_));
 sky130_fd_sc_hd__a221o_1 _11584_ (.A1(\core.count_instr[57] ),
    .A2(_05350_),
    .B1(_05384_),
    .B2(\core.count_cycle[25] ),
    .C1(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__nor2_1 _11585_ (.A(\core.reg_pc[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_2 _11586_ (.A(\core.reg_pc[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_05453_));
 sky130_fd_sc_hd__inv_2 _11587_ (.A(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__nor2_1 _11588_ (.A(_05452_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__inv_2 _11589_ (.A(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_2 _11590_ (.A(_05445_),
    .B(_05433_),
    .Y(_05457_));
 sky130_fd_sc_hd__xor2_1 _11591_ (.A(_05456_),
    .B(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__a21oi_1 _11592_ (.A1(_05317_),
    .A2(net18),
    .B1(_05364_),
    .Y(_05459_));
 sky130_fd_sc_hd__o32a_1 _11593_ (.A1(_05316_),
    .A2(_05459_),
    .A3(_05366_),
    .B1(_05319_),
    .B2(_04942_),
    .X(_05460_));
 sky130_fd_sc_hd__o21ai_1 _11594_ (.A1(_05354_),
    .A2(_05458_),
    .B1(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a21o_1 _11595_ (.A1(_05398_),
    .A2(_05451_),
    .B1(_05461_),
    .X(_01560_));
 sky130_fd_sc_hd__a22o_1 _11596_ (.A1(\core.count_instr[26] ),
    .A2(_05351_),
    .B1(_05385_),
    .B2(\core.count_cycle[58] ),
    .X(_05462_));
 sky130_fd_sc_hd__a221o_1 _11597_ (.A1(\core.count_instr[58] ),
    .A2(_05350_),
    .B1(_05384_),
    .B2(\core.count_cycle[26] ),
    .C1(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_2 _11598_ (.A(\core.reg_pc[26] ),
    .X(_05464_));
 sky130_fd_sc_hd__nor2_1 _11599_ (.A(_05464_),
    .B(\core.decoded_imm[26] ),
    .Y(_05465_));
 sky130_fd_sc_hd__nand2_2 _11600_ (.A(_05464_),
    .B(\core.decoded_imm[26] ),
    .Y(_05466_));
 sky130_fd_sc_hd__and2b_1 _11601_ (.A_N(_05465_),
    .B(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__and2_2 _11602_ (.A(_05435_),
    .B(_05455_),
    .X(_05468_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_05443_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__o21a_1 _11604_ (.A1(_05433_),
    .A2(_05452_),
    .B1(_05453_),
    .X(_05470_));
 sky130_fd_sc_hd__nand2_1 _11605_ (.A(_05469_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__or2_4 _11606_ (.A(_05467_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__nand2_1 _11607_ (.A(_05471_),
    .B(_05467_),
    .Y(_05473_));
 sky130_fd_sc_hd__nand2_2 _11608_ (.A(_05472_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a21oi_1 _11609_ (.A1(_05317_),
    .A2(net19),
    .B1(_05364_),
    .Y(_05475_));
 sky130_fd_sc_hd__o32a_1 _11610_ (.A1(_05316_),
    .A2(_05475_),
    .A3(_05366_),
    .B1(_05319_),
    .B2(_04819_),
    .X(_05476_));
 sky130_fd_sc_hd__o21ai_2 _11611_ (.A1(_05354_),
    .A2(_05474_),
    .B1(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__a21o_1 _11612_ (.A1(_05398_),
    .A2(_05463_),
    .B1(_05477_),
    .X(_01561_));
 sky130_fd_sc_hd__nor2_1 _11613_ (.A(\core.reg_pc[27] ),
    .B(\core.decoded_imm[27] ),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_1 _11614_ (.A(\core.reg_pc[27] ),
    .B(\core.decoded_imm[27] ),
    .Y(_05479_));
 sky130_fd_sc_hd__and2b_2 _11615_ (.A_N(_05478_),
    .B(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__nand2_1 _11616_ (.A(_05473_),
    .B(_05466_),
    .Y(_05481_));
 sky130_fd_sc_hd__or2_1 _11617_ (.A(_05480_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__nand2_2 _11618_ (.A(_05481_),
    .B(_05480_),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_1 _11619_ (.A(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__a21oi_1 _11620_ (.A1(_05363_),
    .A2(net20),
    .B1(_05286_),
    .Y(_05485_));
 sky130_fd_sc_hd__o32a_1 _11621_ (.A1(_05362_),
    .A2(_05485_),
    .A3(_05292_),
    .B1(_05080_),
    .B2(_04814_),
    .X(_05486_));
 sky130_fd_sc_hd__a22o_1 _11622_ (.A1(\core.count_instr[27] ),
    .A2(_05088_),
    .B1(_05296_),
    .B2(\core.count_cycle[59] ),
    .X(_05487_));
 sky130_fd_sc_hd__a221o_1 _11623_ (.A1(\core.count_instr[59] ),
    .A2(_05104_),
    .B1(_05105_),
    .B2(\core.count_cycle[27] ),
    .C1(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__nand2_4 _11624_ (.A(_05488_),
    .B(_05268_),
    .Y(_05489_));
 sky130_fd_sc_hd__o211ai_2 _11625_ (.A1(_04493_),
    .A2(_05484_),
    .B1(_05486_),
    .C1(_05489_),
    .Y(_01562_));
 sky130_fd_sc_hd__a22o_1 _11626_ (.A1(\core.count_instr[28] ),
    .A2(_05295_),
    .B1(_05385_),
    .B2(\core.count_cycle[60] ),
    .X(_05490_));
 sky130_fd_sc_hd__a221o_1 _11627_ (.A1(\core.count_instr[60] ),
    .A2(_05294_),
    .B1(_05384_),
    .B2(\core.count_cycle[28] ),
    .C1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__buf_2 _11628_ (.A(\core.reg_pc[28] ),
    .X(_05492_));
 sky130_fd_sc_hd__nor2_2 _11629_ (.A(_05492_),
    .B(\core.decoded_imm[28] ),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _11630_ (.A(_05492_),
    .B(\core.decoded_imm[28] ),
    .Y(_05494_));
 sky130_fd_sc_hd__and2b_1 _11631_ (.A_N(_05493_),
    .B(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__nand2_1 _11632_ (.A(_05467_),
    .B(_05480_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand3b_1 _11633_ (.A_N(_05496_),
    .B(_05443_),
    .C(_05468_),
    .Y(_05497_));
 sky130_fd_sc_hd__o221a_1 _11634_ (.A1(_05466_),
    .A2(_05478_),
    .B1(_05496_),
    .B2(_05470_),
    .C1(_05479_),
    .X(_05498_));
 sky130_fd_sc_hd__nand2_1 _11635_ (.A(_05497_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__or2_1 _11636_ (.A(_05495_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__nand2_2 _11637_ (.A(_05499_),
    .B(_05495_),
    .Y(_05501_));
 sky130_fd_sc_hd__nand2_2 _11638_ (.A(_05500_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__a21oi_1 _11639_ (.A1(_05317_),
    .A2(net21),
    .B1(_05364_),
    .Y(_05503_));
 sky130_fd_sc_hd__o32a_1 _11640_ (.A1(_05316_),
    .A2(_05503_),
    .A3(_05366_),
    .B1(_05319_),
    .B2(_04931_),
    .X(_05504_));
 sky130_fd_sc_hd__o21ai_1 _11641_ (.A1(_05354_),
    .A2(_05502_),
    .B1(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__a21o_1 _11642_ (.A1(_05398_),
    .A2(_05491_),
    .B1(_05505_),
    .X(_01563_));
 sky130_fd_sc_hd__nor2_1 _11643_ (.A(\core.reg_pc[29] ),
    .B(\core.decoded_imm[29] ),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2_1 _11644_ (.A(\core.reg_pc[29] ),
    .B(\core.decoded_imm[29] ),
    .Y(_05507_));
 sky130_fd_sc_hd__and2b_1 _11645_ (.A_N(_05506_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__nand2_1 _11646_ (.A(_05501_),
    .B(_05494_),
    .Y(_05509_));
 sky130_fd_sc_hd__or2_1 _11647_ (.A(_05508_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__nand2_1 _11648_ (.A(_05509_),
    .B(_05508_),
    .Y(_05511_));
 sky130_fd_sc_hd__nand3_1 _11649_ (.A(_05510_),
    .B(_04982_),
    .C(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__a21oi_1 _11650_ (.A1(_05363_),
    .A2(net22),
    .B1(_05286_),
    .Y(_05513_));
 sky130_fd_sc_hd__o32a_1 _11651_ (.A1(_05362_),
    .A2(_05513_),
    .A3(_05292_),
    .B1(_04587_),
    .B2(_04933_),
    .X(_05514_));
 sky130_fd_sc_hd__a22o_1 _11652_ (.A1(\core.count_instr[29] ),
    .A2(_05295_),
    .B1(_05296_),
    .B2(\core.count_cycle[61] ),
    .X(_05515_));
 sky130_fd_sc_hd__a221o_1 _11653_ (.A1(\core.count_instr[61] ),
    .A2(_05294_),
    .B1(_05037_),
    .B2(\core.count_cycle[29] ),
    .C1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_1 _11654_ (.A(_05516_),
    .B(_05268_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand3_1 _11655_ (.A(_05512_),
    .B(_05514_),
    .C(_05517_),
    .Y(_01564_));
 sky130_fd_sc_hd__inv_2 _11656_ (.A(\core.reg_pc[30] ),
    .Y(_05518_));
 sky130_fd_sc_hd__inv_2 _11657_ (.A(\core.decoded_imm[30] ),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _11658_ (.A(_05518_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_1 _11659_ (.A(\core.reg_pc[30] ),
    .B(\core.decoded_imm[30] ),
    .Y(_05521_));
 sky130_fd_sc_hd__and2_1 _11660_ (.A(_05520_),
    .B(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__and2_1 _11661_ (.A(_05495_),
    .B(_05508_),
    .X(_05523_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_05499_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21a_1 _11663_ (.A1(_05494_),
    .A2(_05506_),
    .B1(_05507_),
    .X(_05525_));
 sky130_fd_sc_hd__nand2_1 _11664_ (.A(_05524_),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__or2_1 _11665_ (.A(_05522_),
    .B(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__nand2_1 _11666_ (.A(_05526_),
    .B(_05522_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand3_1 _11667_ (.A(_05527_),
    .B(_04982_),
    .C(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__a22o_1 _11668_ (.A1(\core.count_instr[30] ),
    .A2(_05295_),
    .B1(_05296_),
    .B2(\core.count_cycle[62] ),
    .X(_05530_));
 sky130_fd_sc_hd__a221o_4 _11669_ (.A1(\core.count_instr[62] ),
    .A2(_05294_),
    .B1(_05037_),
    .B2(\core.count_cycle[30] ),
    .C1(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_05531_),
    .B(_05268_),
    .Y(_05532_));
 sky130_fd_sc_hd__a21oi_1 _11671_ (.A1(_05424_),
    .A2(net24),
    .B1(_05286_),
    .Y(_05533_));
 sky130_fd_sc_hd__o32a_1 _11672_ (.A1(_05068_),
    .A2(_05533_),
    .A3(_05292_),
    .B1(_04587_),
    .B2(_04843_),
    .X(_05534_));
 sky130_fd_sc_hd__nand3_1 _11673_ (.A(_05529_),
    .B(_05532_),
    .C(_05534_),
    .Y(_01566_));
 sky130_fd_sc_hd__nand2_1 _11674_ (.A(_05528_),
    .B(_05521_),
    .Y(_05535_));
 sky130_fd_sc_hd__xor2_1 _11675_ (.A(\core.reg_pc[31] ),
    .B(\core.decoded_imm[31] ),
    .X(_05536_));
 sky130_fd_sc_hd__nand2_1 _11676_ (.A(_05535_),
    .B(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__inv_2 _11677_ (.A(_05536_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand3_2 _11678_ (.A(_05528_),
    .B(_05521_),
    .C(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand3_1 _11679_ (.A(_05537_),
    .B(_04982_),
    .C(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__a21oi_1 _11680_ (.A1(_05363_),
    .A2(net25),
    .B1(_05286_),
    .Y(_05541_));
 sky130_fd_sc_hd__o32a_4 _11681_ (.A1(_05362_),
    .A2(_05541_),
    .A3(_05292_),
    .B1(_04587_),
    .B2(_04838_),
    .X(_05542_));
 sky130_fd_sc_hd__a22o_1 _11682_ (.A1(\core.count_instr[31] ),
    .A2(_05295_),
    .B1(_05296_),
    .B2(\core.count_cycle[63] ),
    .X(_05543_));
 sky130_fd_sc_hd__a221o_2 _11683_ (.A1(\core.count_instr[63] ),
    .A2(_05294_),
    .B1(_05037_),
    .B2(\core.count_cycle[31] ),
    .C1(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__nand2_2 _11684_ (.A(_05544_),
    .B(_05268_),
    .Y(_05545_));
 sky130_fd_sc_hd__nand3_1 _11685_ (.A(_05540_),
    .B(_05542_),
    .C(_05545_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_4 _11686_ (.A(\core.instr_andi ),
    .B(\core.instr_and ),
    .Y(_05546_));
 sky130_fd_sc_hd__inv_2 _11687_ (.A(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__nor2_1 _11688_ (.A(\core.instr_or ),
    .B(\core.instr_ori ),
    .Y(_05548_));
 sky130_fd_sc_hd__inv_2 _11689_ (.A(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__nor2_1 _11690_ (.A(\core.instr_xori ),
    .B(\core.instr_xor ),
    .Y(_05550_));
 sky130_fd_sc_hd__or4b_4 _11691_ (.A(\core.is_compare ),
    .B(_05547_),
    .C(_05549_),
    .D_N(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__clkbuf_2 _11692_ (.A(_05546_),
    .X(_05552_));
 sky130_fd_sc_hd__buf_1 _11693_ (.A(_05548_),
    .X(_05553_));
 sky130_fd_sc_hd__o22a_1 _11694_ (.A1(_04960_),
    .A2(_05552_),
    .B1(_04959_),
    .B2(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__clkbuf_4 _11695_ (.A(_05550_),
    .X(_05555_));
 sky130_fd_sc_hd__or2_1 _11696_ (.A(_05555_),
    .B(_04962_),
    .X(_05556_));
 sky130_fd_sc_hd__nand2_1 _11697_ (.A(_04974_),
    .B(net176),
    .Y(_05557_));
 sky130_fd_sc_hd__o2111ai_1 _11698_ (.A1(_04962_),
    .A2(_05551_),
    .B1(_05554_),
    .C1(_05556_),
    .D1(_05557_),
    .Y(\core.alu_out[0] ));
 sky130_fd_sc_hd__clkinv_4 _11699_ (.A(_05551_),
    .Y(_05558_));
 sky130_fd_sc_hd__buf_2 _11700_ (.A(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__xor2_1 _11701_ (.A(_04695_),
    .B(_04692_),
    .X(_05560_));
 sky130_fd_sc_hd__xor2_1 _11702_ (.A(_04960_),
    .B(_04692_),
    .X(_05561_));
 sky130_fd_sc_hd__inv_2 _11703_ (.A(\core.instr_sub ),
    .Y(_05562_));
 sky130_fd_sc_hd__buf_2 _11704_ (.A(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_4 _11705_ (.A(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11706_ (.A(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(_05560_),
    .A1(_05561_),
    .S(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_8 _11708_ (.A(_05555_),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_4 _11709_ (.A(_05567_),
    .B(_04692_),
    .Y(_05568_));
 sky130_fd_sc_hd__clkbuf_4 _11710_ (.A(_05549_),
    .X(_05569_));
 sky130_fd_sc_hd__a2bb2o_1 _11711_ (.A1_N(_04691_),
    .A2_N(_05546_),
    .B1(_04690_),
    .B2(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__a211o_1 _11712_ (.A1(_05559_),
    .A2(_05566_),
    .B1(_05568_),
    .C1(_05570_),
    .X(\core.alu_out[1] ));
 sky130_fd_sc_hd__inv_2 _11713_ (.A(_04686_),
    .Y(_05571_));
 sky130_fd_sc_hd__clkbuf_4 _11714_ (.A(\core.instr_sub ),
    .X(_05572_));
 sky130_fd_sc_hd__nor2_1 _11715_ (.A(\core.pcpi_rs1[1] ),
    .B(_04696_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21a_1 _11716_ (.A1(_04960_),
    .A2(_05573_),
    .B1(_04691_),
    .X(_05574_));
 sky130_fd_sc_hd__nand2_1 _11717_ (.A(_04698_),
    .B(_05572_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_2 _11718_ (.A1(_05572_),
    .A2(_05574_),
    .B1(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__or2_1 _11719_ (.A(_05571_),
    .B(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_4 _11720_ (.A(_05576_),
    .B(_05571_),
    .Y(_05578_));
 sky130_fd_sc_hd__buf_4 _11721_ (.A(_05550_),
    .X(_05579_));
 sky130_fd_sc_hd__nor2_4 _11722_ (.A(_05579_),
    .B(_04686_),
    .Y(_05580_));
 sky130_fd_sc_hd__a2bb2o_1 _11723_ (.A1_N(_04685_),
    .A2_N(_05546_),
    .B1(_04684_),
    .B2(_05569_),
    .X(_05581_));
 sky130_fd_sc_hd__a311o_1 _11724_ (.A1(_05559_),
    .A2(_05577_),
    .A3(_05578_),
    .B1(_05580_),
    .C1(_05581_),
    .X(\core.alu_out[2] ));
 sky130_fd_sc_hd__o21ai_2 _11725_ (.A1(_04686_),
    .A2(_05574_),
    .B1(_04685_),
    .Y(_05582_));
 sky130_fd_sc_hd__or2_1 _11726_ (.A(_05571_),
    .B(_04698_),
    .X(_05583_));
 sky130_fd_sc_hd__a21oi_1 _11727_ (.A1(_04682_),
    .A2(_04699_),
    .B1(_05562_),
    .Y(_05584_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(_05582_),
    .A2(_05563_),
    .B1(_05583_),
    .B2(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__inv_2 _11729_ (.A(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__or2_2 _11730_ (.A(_04681_),
    .B(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__nand2_2 _11731_ (.A(_05586_),
    .B(_04681_),
    .Y(_05588_));
 sky130_fd_sc_hd__buf_1 _11732_ (.A(_05558_),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_4 _11733_ (.A(_05555_),
    .X(_05590_));
 sky130_fd_sc_hd__nor2_1 _11734_ (.A(_05590_),
    .B(_04681_),
    .Y(_05591_));
 sky130_fd_sc_hd__buf_2 _11735_ (.A(_05547_),
    .X(_05592_));
 sky130_fd_sc_hd__inv_2 _11736_ (.A(_04680_),
    .Y(_05593_));
 sky130_fd_sc_hd__a22o_1 _11737_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_04678_),
    .B2(_05569_),
    .X(_05594_));
 sky130_fd_sc_hd__a311o_1 _11738_ (.A1(_05587_),
    .A2(_05588_),
    .A3(_05589_),
    .B1(_05591_),
    .C1(_05594_),
    .X(\core.alu_out[3] ));
 sky130_fd_sc_hd__inv_2 _11739_ (.A(_04725_),
    .Y(_05595_));
 sky130_fd_sc_hd__buf_2 _11740_ (.A(_05563_),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_2 _11741_ (.A(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__a21o_1 _11742_ (.A1(_05582_),
    .A2(_04678_),
    .B1(_05593_),
    .X(_05598_));
 sky130_fd_sc_hd__clkbuf_2 _11743_ (.A(_05564_),
    .X(_05599_));
 sky130_fd_sc_hd__nand2_1 _11744_ (.A(_05598_),
    .B(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21ai_2 _11745_ (.A1(_05597_),
    .A2(_04703_),
    .B1(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__or2_1 _11746_ (.A(_05595_),
    .B(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__buf_2 _11747_ (.A(_05589_),
    .X(_05603_));
 sky130_fd_sc_hd__nand2_1 _11748_ (.A(_05601_),
    .B(_05595_),
    .Y(_05604_));
 sky130_fd_sc_hd__inv_2 _11749_ (.A(_04724_),
    .Y(_05605_));
 sky130_fd_sc_hd__nor2_1 _11750_ (.A(_05555_),
    .B(_04725_),
    .Y(_05606_));
 sky130_fd_sc_hd__a221o_1 _11751_ (.A1(_04721_),
    .A2(_05549_),
    .B1(_05605_),
    .B2(_05592_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__a31o_1 _11752_ (.A1(_05602_),
    .A2(_05603_),
    .A3(_05604_),
    .B1(_05607_),
    .X(\core.alu_out[4] ));
 sky130_fd_sc_hd__clkbuf_4 _11753_ (.A(\core.instr_sub ),
    .X(_05608_));
 sky130_fd_sc_hd__a21oi_1 _11754_ (.A1(_05598_),
    .A2(_04721_),
    .B1(_05605_),
    .Y(_05609_));
 sky130_fd_sc_hd__a211o_1 _11755_ (.A1(_04703_),
    .A2(_04725_),
    .B1(_05563_),
    .C1(_04731_),
    .X(_05610_));
 sky130_fd_sc_hd__o21ai_2 _11756_ (.A1(_05608_),
    .A2(_05609_),
    .B1(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__or2_1 _11757_ (.A(_04718_),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_4 _11758_ (.A(_05611_),
    .B(_04718_),
    .Y(_05613_));
 sky130_fd_sc_hd__nor2_4 _11759_ (.A(_05590_),
    .B(_04719_),
    .Y(_05614_));
 sky130_fd_sc_hd__a2bb2o_1 _11760_ (.A1_N(_04715_),
    .A2_N(_05548_),
    .B1(_04717_),
    .B2(_05592_),
    .X(_05615_));
 sky130_fd_sc_hd__a311o_1 _11761_ (.A1(_05612_),
    .A2(_05613_),
    .A3(_05589_),
    .B1(_05614_),
    .C1(_05615_),
    .X(\core.alu_out[5] ));
 sky130_fd_sc_hd__inv_2 _11762_ (.A(_04711_),
    .Y(_05616_));
 sky130_fd_sc_hd__clkbuf_2 _11763_ (.A(_05596_),
    .X(_05617_));
 sky130_fd_sc_hd__a31o_1 _11764_ (.A1(_04703_),
    .A2(_04719_),
    .A3(_04725_),
    .B1(_04733_),
    .X(_05618_));
 sky130_fd_sc_hd__nor2_1 _11765_ (.A(_04725_),
    .B(_04719_),
    .Y(_05619_));
 sky130_fd_sc_hd__o21ai_2 _11766_ (.A1(_04724_),
    .A2(_04715_),
    .B1(_04716_),
    .Y(_05620_));
 sky130_fd_sc_hd__a21o_2 _11767_ (.A1(_05598_),
    .A2(_05619_),
    .B1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__nand2_1 _11768_ (.A(_05621_),
    .B(_05599_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_1 _11769_ (.A1(_05617_),
    .A2(_05618_),
    .B1(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__or2_1 _11770_ (.A(_05616_),
    .B(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__nand2_1 _11771_ (.A(_05623_),
    .B(_05616_),
    .Y(_05625_));
 sky130_fd_sc_hd__clkbuf_2 _11772_ (.A(_05546_),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_2 _11773_ (.A(_05555_),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_2 _11774_ (.A(_05549_),
    .X(_05628_));
 sky130_fd_sc_hd__nand2_2 _11775_ (.A(_04708_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__o221ai_1 _11776_ (.A1(_04710_),
    .A2(_05626_),
    .B1(_05627_),
    .B2(_04711_),
    .C1(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__a31o_1 _11777_ (.A1(_05624_),
    .A2(_05603_),
    .A3(_05625_),
    .B1(_05630_),
    .X(\core.alu_out[6] ));
 sky130_fd_sc_hd__clkbuf_4 _11778_ (.A(_05563_),
    .X(_05631_));
 sky130_fd_sc_hd__nand2_2 _11779_ (.A(_05621_),
    .B(_05616_),
    .Y(_05632_));
 sky130_fd_sc_hd__a21o_1 _11780_ (.A1(_05618_),
    .A2(_04711_),
    .B1(_04739_),
    .X(_05633_));
 sky130_fd_sc_hd__and2_1 _11781_ (.A(_05633_),
    .B(\core.instr_sub ),
    .X(_05634_));
 sky130_fd_sc_hd__a31o_1 _11782_ (.A1(_05631_),
    .A2(_04710_),
    .A3(_05632_),
    .B1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__or2_1 _11783_ (.A(_04736_),
    .B(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__nand2_1 _11784_ (.A(_05635_),
    .B(_04736_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_04704_),
    .B(_05628_),
    .Y(_05638_));
 sky130_fd_sc_hd__o221ai_2 _11786_ (.A1(_04706_),
    .A2(_05626_),
    .B1(_05627_),
    .B2(_04736_),
    .C1(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a31o_1 _11787_ (.A1(_05636_),
    .A2(_05603_),
    .A3(_05637_),
    .B1(_05639_),
    .X(\core.alu_out[7] ));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(_04736_),
    .B(_04711_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand3_2 _11789_ (.A(_05598_),
    .B(_05619_),
    .C(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__nand2_4 _11790_ (.A(_05640_),
    .B(_05620_),
    .Y(_05642_));
 sky130_fd_sc_hd__o211a_4 _11791_ (.A1(_04736_),
    .A2(_04710_),
    .B1(_04706_),
    .C1(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_4 _11792_ (.A(_05641_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_05644_),
    .B(_05565_),
    .Y(_05645_));
 sky130_fd_sc_hd__or2_1 _11794_ (.A(_05563_),
    .B(_04743_),
    .X(_05646_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11795_ (.A(_04761_),
    .X(_05647_));
 sky130_fd_sc_hd__a21oi_1 _11796_ (.A1(_05645_),
    .A2(_05646_),
    .B1(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__and3_1 _11797_ (.A(_05645_),
    .B(_05647_),
    .C(_05646_),
    .X(_05649_));
 sky130_fd_sc_hd__or2_1 _11798_ (.A(_04758_),
    .B(_05553_),
    .X(_05650_));
 sky130_fd_sc_hd__o221a_1 _11799_ (.A1(_04759_),
    .A2(_05552_),
    .B1(_05590_),
    .B2(_05647_),
    .C1(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__o31ai_1 _11800_ (.A1(_05551_),
    .A2(_05648_),
    .A3(_05649_),
    .B1(_05651_),
    .Y(\core.alu_out[8] ));
 sky130_fd_sc_hd__a21oi_1 _11801_ (.A1(_04743_),
    .A2(_05647_),
    .B1(_04784_),
    .Y(_05652_));
 sky130_fd_sc_hd__inv_2 _11802_ (.A(_05647_),
    .Y(_05653_));
 sky130_fd_sc_hd__a211o_1 _11803_ (.A1(_05644_),
    .A2(_05653_),
    .B1(\core.instr_sub ),
    .C1(_04760_),
    .X(_05654_));
 sky130_fd_sc_hd__o21ai_2 _11804_ (.A1(_05617_),
    .A2(_05652_),
    .B1(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(_04757_),
    .B(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__nand2_2 _11806_ (.A(_05655_),
    .B(_04757_),
    .Y(_05657_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11807_ (.A(_05548_),
    .X(_05658_));
 sky130_fd_sc_hd__buf_2 _11808_ (.A(_05547_),
    .X(_05659_));
 sky130_fd_sc_hd__nand2_2 _11809_ (.A(_05659_),
    .B(_04755_),
    .Y(_05660_));
 sky130_fd_sc_hd__o221ai_1 _11810_ (.A1(_04753_),
    .A2(_05658_),
    .B1(_05627_),
    .B2(_04757_),
    .C1(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__a31o_1 _11811_ (.A1(_05656_),
    .A2(_05603_),
    .A3(_05657_),
    .B1(_05661_),
    .X(\core.alu_out[9] ));
 sky130_fd_sc_hd__inv_2 _11812_ (.A(_04750_),
    .Y(_05662_));
 sky130_fd_sc_hd__and2_1 _11813_ (.A(_04727_),
    .B(_04742_),
    .X(_05663_));
 sky130_fd_sc_hd__o211a_1 _11814_ (.A1(_04762_),
    .A2(_05663_),
    .B1(_04787_),
    .C1(_04785_),
    .X(_05664_));
 sky130_fd_sc_hd__nor2_1 _11815_ (.A(_04757_),
    .B(_05647_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_2 _11816_ (.A1(_04759_),
    .A2(_04753_),
    .B1(_04754_),
    .Y(_05666_));
 sky130_fd_sc_hd__a21o_1 _11817_ (.A1(_05644_),
    .A2(_05665_),
    .B1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(_05664_),
    .A1(_05667_),
    .S(_05564_),
    .X(_05668_));
 sky130_fd_sc_hd__or2_1 _11819_ (.A(_05662_),
    .B(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_2 _11820_ (.A(_05668_),
    .B(_05662_),
    .Y(_05670_));
 sky130_fd_sc_hd__nand2_1 _11821_ (.A(_04748_),
    .B(_05628_),
    .Y(_05671_));
 sky130_fd_sc_hd__o221ai_1 _11822_ (.A1(_04749_),
    .A2(_05626_),
    .B1(_05627_),
    .B2(_04750_),
    .C1(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__a31o_1 _11823_ (.A1(_05669_),
    .A2(_05603_),
    .A3(_05670_),
    .B1(_05672_),
    .X(\core.alu_out[10] ));
 sky130_fd_sc_hd__nor2_1 _11824_ (.A(_05662_),
    .B(_05664_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21ai_1 _11825_ (.A1(_04791_),
    .A2(_05673_),
    .B1(_05608_),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _11826_ (.A(_04749_),
    .B(_05564_),
    .Y(_05675_));
 sky130_fd_sc_hd__a21o_1 _11827_ (.A1(_05667_),
    .A2(_05662_),
    .B1(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_05674_),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__or2_1 _11829_ (.A(_04789_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_2 _11830_ (.A(_05558_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(_05677_),
    .B(_04789_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand2_4 _11832_ (.A(_05659_),
    .B(_04746_),
    .Y(_05681_));
 sky130_fd_sc_hd__o221ai_2 _11833_ (.A1(_04744_),
    .A2(_05658_),
    .B1(_05627_),
    .B2(_04789_),
    .C1(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a31o_1 _11834_ (.A1(_05678_),
    .A2(_05679_),
    .A3(_05680_),
    .B1(_05682_),
    .X(\core.alu_out[11] ));
 sky130_fd_sc_hd__inv_2 _11835_ (.A(_04778_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _11836_ (.A(_04743_),
    .B(_04763_),
    .Y(_05684_));
 sky130_fd_sc_hd__inv_2 _11837_ (.A(_04795_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_2 _11838_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__nor2_1 _11839_ (.A(_04750_),
    .B(_04789_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(_05665_),
    .B(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__inv_2 _11841_ (.A(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__nor2_1 _11842_ (.A(_04749_),
    .B(_04789_),
    .Y(_05690_));
 sky130_fd_sc_hd__a211o_1 _11843_ (.A1(_05687_),
    .A2(_05666_),
    .B1(_04746_),
    .C1(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__a21o_1 _11844_ (.A1(_05644_),
    .A2(_05689_),
    .B1(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_05692_),
    .B(_05631_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_2 _11846_ (.A1(_05631_),
    .A2(_05686_),
    .B1(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__or2_1 _11847_ (.A(_05683_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_4 _11848_ (.A(_05694_),
    .B(_05683_),
    .Y(_05696_));
 sky130_fd_sc_hd__nor2_4 _11849_ (.A(_05590_),
    .B(_04778_),
    .Y(_05697_));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(_04777_),
    .Y(_05698_));
 sky130_fd_sc_hd__a22o_1 _11851_ (.A1(_05592_),
    .A2(_05698_),
    .B1(_04776_),
    .B2(_05569_),
    .X(_05699_));
 sky130_fd_sc_hd__a311o_1 _11852_ (.A1(_05695_),
    .A2(_05696_),
    .A3(_05589_),
    .B1(_05697_),
    .C1(_05699_),
    .X(\core.alu_out[12] ));
 sky130_fd_sc_hd__a21o_1 _11853_ (.A1(_05686_),
    .A2(_04778_),
    .B1(_04797_),
    .X(_05700_));
 sky130_fd_sc_hd__nand2_4 _11854_ (.A(_05692_),
    .B(_05683_),
    .Y(_05701_));
 sky130_fd_sc_hd__nor2_1 _11855_ (.A(_05572_),
    .B(_05698_),
    .Y(_05702_));
 sky130_fd_sc_hd__a22o_1 _11856_ (.A1(_05700_),
    .A2(_05572_),
    .B1(_05701_),
    .B2(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__or2_1 _11857_ (.A(_04775_),
    .B(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__nand2_1 _11858_ (.A(_05703_),
    .B(_04775_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_4 _11859_ (.A(_05659_),
    .B(_04773_),
    .Y(_05706_));
 sky130_fd_sc_hd__o221ai_1 _11860_ (.A1(_04771_),
    .A2(_05658_),
    .B1(_05627_),
    .B2(_04775_),
    .C1(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__a31o_1 _11861_ (.A1(_05704_),
    .A2(_05679_),
    .A3(_05705_),
    .B1(_05707_),
    .X(\core.alu_out[13] ));
 sky130_fd_sc_hd__inv_2 _11862_ (.A(_05686_),
    .Y(_05708_));
 sky130_fd_sc_hd__o21a_1 _11863_ (.A1(_04779_),
    .A2(_05708_),
    .B1(_04802_),
    .X(_05709_));
 sky130_fd_sc_hd__nor2_1 _11864_ (.A(_04778_),
    .B(_04775_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21a_1 _11865_ (.A1(_04777_),
    .A2(_04771_),
    .B1(_04772_),
    .X(_05711_));
 sky130_fd_sc_hd__inv_2 _11866_ (.A(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__a21oi_1 _11867_ (.A1(_05692_),
    .A2(_05710_),
    .B1(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _11868_ (.A(_05713_),
    .B(_05599_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_2 _11869_ (.A1(_05617_),
    .A2(_05709_),
    .B1(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__or2_1 _11870_ (.A(_04769_),
    .B(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__nand2_2 _11871_ (.A(_05715_),
    .B(_04769_),
    .Y(_05717_));
 sky130_fd_sc_hd__buf_2 _11872_ (.A(_05555_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_2 _11873_ (.A(_04767_),
    .B(_05628_),
    .Y(_05719_));
 sky130_fd_sc_hd__o221ai_1 _11874_ (.A1(_04768_),
    .A2(_05626_),
    .B1(_05718_),
    .B2(_04769_),
    .C1(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__a31o_1 _11875_ (.A1(_05716_),
    .A2(_05679_),
    .A3(_05717_),
    .B1(_05720_),
    .X(\core.alu_out[14] ));
 sky130_fd_sc_hd__o211ai_2 _11876_ (.A1(_04769_),
    .A2(_05713_),
    .B1(_05599_),
    .C1(_04768_),
    .Y(_05721_));
 sky130_fd_sc_hd__a21oi_1 _11877_ (.A1(_04767_),
    .A2(_04768_),
    .B1(_05709_),
    .Y(_05722_));
 sky130_fd_sc_hd__o21ai_1 _11878_ (.A1(_04805_),
    .A2(_05722_),
    .B1(_05608_),
    .Y(_05723_));
 sky130_fd_sc_hd__nand2_1 _11879_ (.A(_05721_),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__or2_1 _11880_ (.A(_04803_),
    .B(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11881_ (.A(_05589_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _11882_ (.A(_05724_),
    .B(_04803_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand3_1 _11883_ (.A(_05725_),
    .B(_05726_),
    .C(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__clkbuf_2 _11884_ (.A(_05546_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_4 _11885_ (.A(_05549_),
    .X(_05730_));
 sky130_fd_sc_hd__nand2_4 _11886_ (.A(_04764_),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__o221a_4 _11887_ (.A1(_04765_),
    .A2(_05729_),
    .B1(_05567_),
    .B2(_04803_),
    .C1(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_1 _11888_ (.A(_05728_),
    .B(_05732_),
    .Y(\core.alu_out[15] ));
 sky130_fd_sc_hd__inv_2 _11889_ (.A(_04873_),
    .Y(_05733_));
 sky130_fd_sc_hd__nor2_1 _11890_ (.A(_04803_),
    .B(_04769_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand2_1 _11891_ (.A(_05710_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__inv_2 _11892_ (.A(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand3_2 _11893_ (.A(_05644_),
    .B(_05689_),
    .C(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21ai_1 _11894_ (.A1(_04768_),
    .A2(_04803_),
    .B1(_04765_),
    .Y(_05738_));
 sky130_fd_sc_hd__a21o_1 _11895_ (.A1(_05712_),
    .A2(_05734_),
    .B1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__a21oi_2 _11896_ (.A1(_05691_),
    .A2(_05736_),
    .B1(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_4 _11897_ (.A(_05737_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _11898_ (.A(_05741_),
    .B(_05596_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21ai_2 _11899_ (.A1(_05631_),
    .A2(_04812_),
    .B1(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__or2_1 _11900_ (.A(_05733_),
    .B(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_4 _11901_ (.A(_05743_),
    .B(_05733_),
    .Y(_05745_));
 sky130_fd_sc_hd__nor2_4 _11902_ (.A(_05590_),
    .B(_04873_),
    .Y(_05746_));
 sky130_fd_sc_hd__inv_2 _11903_ (.A(_04872_),
    .Y(_05747_));
 sky130_fd_sc_hd__a22o_1 _11904_ (.A1(_05592_),
    .A2(_05747_),
    .B1(_04871_),
    .B2(_05569_),
    .X(_05748_));
 sky130_fd_sc_hd__a311o_1 _11905_ (.A1(_05744_),
    .A2(_05745_),
    .A3(_05589_),
    .B1(_05746_),
    .C1(_05748_),
    .X(\core.alu_out[16] ));
 sky130_fd_sc_hd__a21oi_1 _11906_ (.A1(_04812_),
    .A2(_04873_),
    .B1(_04902_),
    .Y(_05749_));
 sky130_fd_sc_hd__a211o_1 _11907_ (.A1(_05741_),
    .A2(_04871_),
    .B1(_05572_),
    .C1(_05747_),
    .X(_05750_));
 sky130_fd_sc_hd__o21ai_1 _11908_ (.A1(_05597_),
    .A2(_05749_),
    .B1(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__or2_1 _11909_ (.A(_04870_),
    .B(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__nand2_1 _11910_ (.A(_05751_),
    .B(_04870_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand3_1 _11911_ (.A(_05752_),
    .B(_05726_),
    .C(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _11912_ (.A(_05659_),
    .B(_04868_),
    .Y(_05755_));
 sky130_fd_sc_hd__o221a_1 _11913_ (.A1(_04866_),
    .A2(_05658_),
    .B1(_05567_),
    .B2(_04870_),
    .C1(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__nand2_1 _11914_ (.A(_05754_),
    .B(_05756_),
    .Y(\core.alu_out[17] ));
 sky130_fd_sc_hd__inv_2 _11915_ (.A(_04876_),
    .Y(_05757_));
 sky130_fd_sc_hd__a31o_1 _11916_ (.A1(_04812_),
    .A2(_04873_),
    .A3(_04870_),
    .B1(_04906_),
    .X(_05758_));
 sky130_fd_sc_hd__o21a_1 _11917_ (.A1(_04872_),
    .A2(_04866_),
    .B1(_04867_),
    .X(_05759_));
 sky130_fd_sc_hd__inv_2 _11918_ (.A(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__a31o_1 _11919_ (.A1(_05741_),
    .A2(_05733_),
    .A3(_04869_),
    .B1(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__nand2_1 _11920_ (.A(_05761_),
    .B(_05631_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_2 _11921_ (.A1(_05631_),
    .A2(_05758_),
    .B1(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nor2_2 _11922_ (.A(_05757_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__and2_1 _11923_ (.A(_05763_),
    .B(_05757_),
    .X(_05765_));
 sky130_fd_sc_hd__nand2_4 _11924_ (.A(_04874_),
    .B(_05569_),
    .Y(_05766_));
 sky130_fd_sc_hd__o221a_1 _11925_ (.A1(_04875_),
    .A2(_05552_),
    .B1(_05590_),
    .B2(_04876_),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__o31ai_2 _11926_ (.A1(_05551_),
    .A2(_05764_),
    .A3(_05765_),
    .B1(_05767_),
    .Y(\core.alu_out[18] ));
 sky130_fd_sc_hd__nand2_1 _11927_ (.A(_04875_),
    .B(_05596_),
    .Y(_05768_));
 sky130_fd_sc_hd__a21o_1 _11928_ (.A1(_05761_),
    .A2(_05757_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__a21o_2 _11929_ (.A1(_05758_),
    .A2(_04876_),
    .B1(_04910_),
    .X(_05770_));
 sky130_fd_sc_hd__nand2_1 _11930_ (.A(_05770_),
    .B(_05608_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _11931_ (.A(_05769_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__or2_1 _11932_ (.A(_04907_),
    .B(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_1 _11933_ (.A(_05772_),
    .B(_04907_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand3_1 _11934_ (.A(_05773_),
    .B(_05726_),
    .C(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_1 _11935_ (.A(_05592_),
    .B(_04864_),
    .Y(_05776_));
 sky130_fd_sc_hd__o221a_1 _11936_ (.A1(_04862_),
    .A2(_05553_),
    .B1(_05579_),
    .B2(_04907_),
    .C1(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__nand2_1 _11937_ (.A(_05775_),
    .B(_05777_),
    .Y(\core.alu_out[19] ));
 sky130_fd_sc_hd__inv_2 _11938_ (.A(_04889_),
    .Y(_05778_));
 sky130_fd_sc_hd__a21o_1 _11939_ (.A1(_04812_),
    .A2(_04877_),
    .B1(_04914_),
    .X(_05779_));
 sky130_fd_sc_hd__nor2_1 _11940_ (.A(_04876_),
    .B(_04907_),
    .Y(_05780_));
 sky130_fd_sc_hd__and3_1 _11941_ (.A(_05780_),
    .B(_05733_),
    .C(_04869_),
    .X(_05781_));
 sky130_fd_sc_hd__nand2_1 _11942_ (.A(_05741_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__nor2_2 _11943_ (.A(_04875_),
    .B(_04907_),
    .Y(_05783_));
 sky130_fd_sc_hd__a211o_1 _11944_ (.A1(_05780_),
    .A2(_05760_),
    .B1(_04864_),
    .C1(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__inv_2 _11945_ (.A(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_2 _11946_ (.A(_05782_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _11947_ (.A(_05786_),
    .B(_05565_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_1 _11948_ (.A1(_05617_),
    .A2(_05779_),
    .B1(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__or2_1 _11949_ (.A(_05778_),
    .B(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _11950_ (.A(_05788_),
    .B(_05778_),
    .Y(_05790_));
 sky130_fd_sc_hd__or2_1 _11951_ (.A(_04886_),
    .B(_05553_),
    .X(_05791_));
 sky130_fd_sc_hd__o221ai_2 _11952_ (.A1(_04887_),
    .A2(_05626_),
    .B1(_05718_),
    .B2(_04889_),
    .C1(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__a31o_1 _11953_ (.A1(_05789_),
    .A2(_05679_),
    .A3(_05790_),
    .B1(_05792_),
    .X(\core.alu_out[20] ));
 sky130_fd_sc_hd__a21oi_1 _11954_ (.A1(_05779_),
    .A2(_04889_),
    .B1(_04918_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_2 _11955_ (.A(_04887_),
    .B(_05564_),
    .Y(_05794_));
 sky130_fd_sc_hd__a21o_1 _11956_ (.A1(_05786_),
    .A2(_05778_),
    .B1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__o21ai_2 _11957_ (.A1(_05617_),
    .A2(_05793_),
    .B1(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__or2_1 _11958_ (.A(_04894_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__nand2_1 _11959_ (.A(_05796_),
    .B(_04894_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _11960_ (.A(_05659_),
    .B(_04892_),
    .Y(_05799_));
 sky130_fd_sc_hd__o221ai_1 _11961_ (.A1(_04890_),
    .A2(_05658_),
    .B1(_05718_),
    .B2(_04894_),
    .C1(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__a31o_1 _11962_ (.A1(_05797_),
    .A2(_05679_),
    .A3(_05798_),
    .B1(_05800_),
    .X(\core.alu_out[21] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11963_ (.A(_04884_),
    .X(_05801_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _11964_ (.A(_05572_),
    .X(_05802_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(_04889_),
    .B(_04894_),
    .Y(_05803_));
 sky130_fd_sc_hd__o21a_1 _11966_ (.A1(_04887_),
    .A2(_04890_),
    .B1(_04891_),
    .X(_05804_));
 sky130_fd_sc_hd__inv_2 _11967_ (.A(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__a21o_1 _11968_ (.A1(_05786_),
    .A2(_05803_),
    .B1(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__a21oi_1 _11969_ (.A1(_04812_),
    .A2(_04877_),
    .B1(_04914_),
    .Y(_05807_));
 sky130_fd_sc_hd__o21bai_2 _11970_ (.A1(_04895_),
    .A2(_05807_),
    .B1_N(_04920_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(_05808_),
    .B(_05802_),
    .Y(_05809_));
 sky130_fd_sc_hd__o21ai_1 _11972_ (.A1(_05802_),
    .A2(_05806_),
    .B1(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__nor2_1 _11973_ (.A(_05801_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__a21o_1 _11974_ (.A1(_05810_),
    .A2(_05801_),
    .B1(_05551_),
    .X(_05812_));
 sky130_fd_sc_hd__nand2_4 _11975_ (.A(_04882_),
    .B(_05730_),
    .Y(_05813_));
 sky130_fd_sc_hd__o221a_1 _11976_ (.A1(_04883_),
    .A2(_05729_),
    .B1(_05567_),
    .B2(_05801_),
    .C1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__o21ai_1 _11977_ (.A1(_05811_),
    .A2(_05812_),
    .B1(_05814_),
    .Y(\core.alu_out[22] ));
 sky130_fd_sc_hd__a21oi_1 _11978_ (.A1(_05786_),
    .A2(_05803_),
    .B1(_05805_),
    .Y(_05815_));
 sky130_fd_sc_hd__o211ai_1 _11979_ (.A1(_05801_),
    .A2(_05815_),
    .B1(_05597_),
    .C1(_04883_),
    .Y(_05816_));
 sky130_fd_sc_hd__a21o_1 _11980_ (.A1(_05808_),
    .A2(_05801_),
    .B1(_04925_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _11981_ (.A(_05817_),
    .B(_05802_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _11982_ (.A(_05816_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(_05819_),
    .B(_04923_),
    .Y(_05820_));
 sky130_fd_sc_hd__nand3b_1 _11984_ (.A_N(_04923_),
    .B(_05816_),
    .C(_05818_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand3_2 _11985_ (.A(_05820_),
    .B(_05821_),
    .C(_05726_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_1 _11986_ (.A(_04878_),
    .B(_05730_),
    .Y(_05823_));
 sky130_fd_sc_hd__o221a_1 _11987_ (.A1(_04880_),
    .A2(_05729_),
    .B1(_05579_),
    .B2(_04923_),
    .C1(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__nand2_1 _11988_ (.A(_05822_),
    .B(_05824_),
    .Y(\core.alu_out[23] ));
 sky130_fd_sc_hd__inv_2 _11989_ (.A(_04811_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21bai_4 _11990_ (.A1(_04897_),
    .A2(_05825_),
    .B1_N(_04929_),
    .Y(_05826_));
 sky130_fd_sc_hd__nor2_2 _11991_ (.A(_05801_),
    .B(_04923_),
    .Y(_05827_));
 sky130_fd_sc_hd__and3_1 _11992_ (.A(_05781_),
    .B(_05803_),
    .C(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__nand2_1 _11993_ (.A(_05741_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_1 _11994_ (.A1(_04883_),
    .A2(_04923_),
    .B1(_04880_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21o_1 _11995_ (.A1(_05805_),
    .A2(_05827_),
    .B1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__a31oi_4 _11996_ (.A1(_05784_),
    .A2(_05803_),
    .A3(_05827_),
    .B1(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_05829_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _11998_ (.A(_05833_),
    .B(_05565_),
    .Y(_05834_));
 sky130_fd_sc_hd__o21ai_1 _11999_ (.A1(_05617_),
    .A2(_05826_),
    .B1(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__or2_1 _12000_ (.A(_04833_),
    .B(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _12001_ (.A(_05835_),
    .B(_04833_),
    .Y(_05837_));
 sky130_fd_sc_hd__or2_1 _12002_ (.A(_04830_),
    .B(_05553_),
    .X(_05838_));
 sky130_fd_sc_hd__o221ai_2 _12003_ (.A1(_04831_),
    .A2(_05626_),
    .B1(_05718_),
    .B2(_04834_),
    .C1(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__a31o_1 _12004_ (.A1(_05836_),
    .A2(_05679_),
    .A3(_05837_),
    .B1(_05839_),
    .X(\core.alu_out[24] ));
 sky130_fd_sc_hd__a21oi_1 _12005_ (.A1(_05826_),
    .A2(_04834_),
    .B1(_04940_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _12006_ (.A(_04831_),
    .B(_05564_),
    .Y(_05841_));
 sky130_fd_sc_hd__a21o_1 _12007_ (.A1(_05833_),
    .A2(_04833_),
    .B1(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__o21ai_2 _12008_ (.A1(_05599_),
    .A2(_05840_),
    .B1(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__or2_1 _12009_ (.A(_04828_),
    .B(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__nand2_1 _12010_ (.A(_05843_),
    .B(_04828_),
    .Y(_05845_));
 sky130_fd_sc_hd__nand2_1 _12011_ (.A(_05659_),
    .B(_04826_),
    .Y(_05846_));
 sky130_fd_sc_hd__o221ai_1 _12012_ (.A1(_04824_),
    .A2(_05658_),
    .B1(_05718_),
    .B2(_04828_),
    .C1(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__a31o_1 _12013_ (.A1(_05844_),
    .A2(_05559_),
    .A3(_05845_),
    .B1(_05847_),
    .X(\core.alu_out[25] ));
 sky130_fd_sc_hd__inv_2 _12014_ (.A(_04822_),
    .Y(_05848_));
 sky130_fd_sc_hd__nor2_1 _12015_ (.A(_04834_),
    .B(_04828_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21a_1 _12016_ (.A1(_04831_),
    .A2(_04824_),
    .B1(_04825_),
    .X(_05850_));
 sky130_fd_sc_hd__a21bo_1 _12017_ (.A1(_05833_),
    .A2(_05849_),
    .B1_N(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__inv_2 _12018_ (.A(_04835_),
    .Y(_05852_));
 sky130_fd_sc_hd__a21oi_2 _12019_ (.A1(_05826_),
    .A2(_05852_),
    .B1(_04944_),
    .Y(_05853_));
 sky130_fd_sc_hd__or2_1 _12020_ (.A(_05596_),
    .B(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__o21a_1 _12021_ (.A1(_05608_),
    .A2(_05851_),
    .B1(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__nor2_1 _12022_ (.A(_05848_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _12023_ (.A(_05855_),
    .B(_05848_),
    .Y(_05857_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(_05857_),
    .B(_05559_),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_05628_),
    .B(_04820_),
    .Y(_05859_));
 sky130_fd_sc_hd__o221a_2 _12026_ (.A1(_04821_),
    .A2(_05729_),
    .B1(_05567_),
    .B2(_04822_),
    .C1(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__o21ai_4 _12027_ (.A1(_05856_),
    .A2(_05858_),
    .B1(_05860_),
    .Y(\core.alu_out[26] ));
 sky130_fd_sc_hd__nand2_2 _12028_ (.A(_04821_),
    .B(_05597_),
    .Y(_05861_));
 sky130_fd_sc_hd__a21o_1 _12029_ (.A1(_05851_),
    .A2(_05848_),
    .B1(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__o21ai_1 _12030_ (.A1(_05848_),
    .A2(_05853_),
    .B1(_04946_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _12031_ (.A(_05863_),
    .B(_05802_),
    .Y(_05864_));
 sky130_fd_sc_hd__nand2_1 _12032_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05865_),
    .B(_04817_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand3_1 _12034_ (.A(_05862_),
    .B(_04947_),
    .C(_05864_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand3_1 _12035_ (.A(_05866_),
    .B(_05726_),
    .C(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nand2_2 _12036_ (.A(_05730_),
    .B(_04815_),
    .Y(_05869_));
 sky130_fd_sc_hd__o221a_1 _12037_ (.A1(_04816_),
    .A2(_05552_),
    .B1(_05579_),
    .B2(_04817_),
    .C1(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__nand2_1 _12038_ (.A(_05868_),
    .B(_05870_),
    .Y(\core.alu_out[27] ));
 sky130_fd_sc_hd__nand2_1 _12039_ (.A(_05826_),
    .B(_04836_),
    .Y(_05871_));
 sky130_fd_sc_hd__inv_2 _12040_ (.A(_04950_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_1 _12041_ (.A(_05871_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__and3_1 _12042_ (.A(_05849_),
    .B(_04947_),
    .C(_05848_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_1 _12043_ (.A(_05833_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_2 _12044_ (.A(_04947_),
    .B(_05848_),
    .Y(_05876_));
 sky130_fd_sc_hd__o221a_4 _12045_ (.A1(_04817_),
    .A2(_04821_),
    .B1(_05850_),
    .B2(_05876_),
    .C1(_04816_),
    .X(_05877_));
 sky130_fd_sc_hd__nand2_2 _12046_ (.A(_05875_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_05878_),
    .B(_05565_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_2 _12048_ (.A1(_05599_),
    .A2(_05873_),
    .B1(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__or2_1 _12049_ (.A(_04853_),
    .B(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_1 _12050_ (.A(_05880_),
    .B(_04853_),
    .Y(_05882_));
 sky130_fd_sc_hd__or2_1 _12051_ (.A(_04850_),
    .B(_05553_),
    .X(_05883_));
 sky130_fd_sc_hd__o221ai_1 _12052_ (.A1(_04851_),
    .A2(_05729_),
    .B1(_05718_),
    .B2(_04854_),
    .C1(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__a31o_1 _12053_ (.A1(_05881_),
    .A2(_05559_),
    .A3(_05882_),
    .B1(_05884_),
    .X(\core.alu_out[28] ));
 sky130_fd_sc_hd__nand2_1 _12054_ (.A(_04851_),
    .B(_05596_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21o_1 _12055_ (.A1(_05878_),
    .A2(_04853_),
    .B1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__a21o_1 _12056_ (.A1(_05873_),
    .A2(_04854_),
    .B1(_04932_),
    .X(_05887_));
 sky130_fd_sc_hd__nand2_1 _12057_ (.A(_05887_),
    .B(_05608_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _12058_ (.A(_05886_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__or2_1 _12059_ (.A(_04930_),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _12060_ (.A(_05889_),
    .B(_04930_),
    .Y(_05891_));
 sky130_fd_sc_hd__nand3_1 _12061_ (.A(_05890_),
    .B(_05726_),
    .C(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__nand2_4 _12062_ (.A(_04855_),
    .B(_05730_),
    .Y(_05893_));
 sky130_fd_sc_hd__o221a_2 _12063_ (.A1(_04857_),
    .A2(_05552_),
    .B1(_05579_),
    .B2(_04930_),
    .C1(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__nand2_4 _12064_ (.A(_05892_),
    .B(_05894_),
    .Y(\core.alu_out[29] ));
 sky130_fd_sc_hd__inv_2 _12065_ (.A(_04847_),
    .Y(_05895_));
 sky130_fd_sc_hd__inv_2 _12066_ (.A(_04859_),
    .Y(_05896_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(_05873_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _12068_ (.A(_05897_),
    .B(_04935_),
    .Y(_05898_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_04930_),
    .B(_04854_),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _12070_ (.A(_05878_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o21a_1 _12071_ (.A1(_04851_),
    .A2(_04930_),
    .B1(_04857_),
    .X(_05901_));
 sky130_fd_sc_hd__nand2_1 _12072_ (.A(_05900_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__nand2_1 _12073_ (.A(_05902_),
    .B(_05597_),
    .Y(_05903_));
 sky130_fd_sc_hd__o21ai_1 _12074_ (.A1(_05597_),
    .A2(_05898_),
    .B1(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__nor2_1 _12075_ (.A(_05895_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_05904_),
    .B(_05895_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_1 _12077_ (.A(_05906_),
    .B(_05559_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_4 _12078_ (.A(_05628_),
    .B(_04844_),
    .Y(_05908_));
 sky130_fd_sc_hd__o221a_1 _12079_ (.A1(_04846_),
    .A2(_05729_),
    .B1(_05567_),
    .B2(_04847_),
    .C1(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__o21ai_1 _12080_ (.A1(_05905_),
    .A2(_05907_),
    .B1(_05909_),
    .Y(\core.alu_out[30] ));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_05898_),
    .B(_04847_),
    .Y(_05910_));
 sky130_fd_sc_hd__o21ai_1 _12082_ (.A1(\core.pcpi_rs2[30] ),
    .A2(_04843_),
    .B1(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_05911_),
    .B(_05802_),
    .Y(_05912_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05902_),
    .B(_05895_),
    .Y(_05913_));
 sky130_fd_sc_hd__and2_1 _12085_ (.A(_04846_),
    .B(_05565_),
    .X(_05914_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_05913_),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__nand2_1 _12087_ (.A(_05912_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _12088_ (.A(_05916_),
    .B(_04841_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand3b_1 _12089_ (.A_N(_04841_),
    .B(_05912_),
    .C(_05915_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand3_1 _12090_ (.A(_05917_),
    .B(_05918_),
    .C(_05603_),
    .Y(_05919_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_05730_),
    .B(_04839_),
    .Y(_05920_));
 sky130_fd_sc_hd__o221a_1 _12092_ (.A1(_04840_),
    .A2(_05552_),
    .B1(_05579_),
    .B2(_04841_),
    .C1(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__nand2_1 _12093_ (.A(_05919_),
    .B(_05921_),
    .Y(\core.alu_out[31] ));
 sky130_fd_sc_hd__clkbuf_2 _12094_ (.A(_04372_),
    .X(_05922_));
 sky130_fd_sc_hd__clkbuf_2 _12095_ (.A(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__clkbuf_2 _12096_ (.A(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(net7),
    .A1(\core.mem_rdata_q[15] ),
    .S(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__clkbuf_1 _12098_ (.A(_05925_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _12099_ (.A0(_01358_),
    .A1(\core.decoded_imm_j[15] ),
    .S(_04979_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _12100_ (.A(_05926_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _12101_ (.A0(net8),
    .A1(\core.mem_rdata_q[16] ),
    .S(_05924_),
    .X(_05927_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12102_ (.A(_05927_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _12103_ (.A0(_01359_),
    .A1(\core.decoded_imm_j[16] ),
    .S(_04979_),
    .X(_05928_));
 sky130_fd_sc_hd__buf_1 _12104_ (.A(_05928_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _12105_ (.A0(net9),
    .A1(\core.mem_rdata_q[17] ),
    .S(_05924_),
    .X(_05929_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12106_ (.A(_05929_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _12107_ (.A0(_01360_),
    .A1(\core.decoded_imm_j[17] ),
    .S(_04979_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_1 _12108_ (.A(_05930_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _12109_ (.A0(net10),
    .A1(\core.mem_rdata_q[18] ),
    .S(_05924_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_2 _12110_ (.A(_05931_),
    .X(_01361_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12111_ (.A(_04977_),
    .X(_05932_));
 sky130_fd_sc_hd__clkbuf_4 _12112_ (.A(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(_01361_),
    .A1(\core.decoded_imm_j[18] ),
    .S(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__clkbuf_8 _12114_ (.A(_05934_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(net11),
    .A1(\core.mem_rdata_q[19] ),
    .S(_05924_),
    .X(_05935_));
 sky130_fd_sc_hd__clkbuf_1 _12116_ (.A(_05935_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(_01362_),
    .A1(\core.decoded_imm_j[19] ),
    .S(_05933_),
    .X(_05936_));
 sky130_fd_sc_hd__buf_1 _12118_ (.A(_05936_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _12119_ (.A0(net13),
    .A1(\core.mem_rdata_q[20] ),
    .S(_05924_),
    .X(_05937_));
 sky130_fd_sc_hd__clkbuf_1 _12120_ (.A(_05937_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _12121_ (.A0(_01363_),
    .A1(_04577_),
    .S(_05933_),
    .X(_05938_));
 sky130_fd_sc_hd__clkbuf_1 _12122_ (.A(_05938_),
    .X(_00020_));
 sky130_fd_sc_hd__clkbuf_2 _12123_ (.A(_05922_),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_2 _12124_ (.A(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(net14),
    .A1(\core.mem_rdata_q[21] ),
    .S(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_2 _12126_ (.A(_05941_),
    .X(_01364_));
 sky130_fd_sc_hd__buf_2 _12127_ (.A(\core.decoded_imm_j[1] ),
    .X(_05942_));
 sky130_fd_sc_hd__mux2_1 _12128_ (.A0(_01364_),
    .A1(_05942_),
    .S(_05933_),
    .X(_05943_));
 sky130_fd_sc_hd__clkbuf_1 _12129_ (.A(_05943_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _12130_ (.A0(net15),
    .A1(\core.mem_rdata_q[22] ),
    .S(_05940_),
    .X(_05944_));
 sky130_fd_sc_hd__clkbuf_2 _12131_ (.A(_05944_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(_01365_),
    .A1(\core.decoded_imm_j[2] ),
    .S(_05933_),
    .X(_05945_));
 sky130_fd_sc_hd__clkbuf_1 _12133_ (.A(_05945_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(net16),
    .A1(\core.mem_rdata_q[23] ),
    .S(_05940_),
    .X(_05946_));
 sky130_fd_sc_hd__buf_1 _12135_ (.A(_05946_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _12136_ (.A0(_01366_),
    .A1(_04575_),
    .S(_05933_),
    .X(_05947_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12137_ (.A(_05947_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(net17),
    .A1(\core.mem_rdata_q[24] ),
    .S(_05940_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_2 _12139_ (.A(_05948_),
    .X(_01367_));
 sky130_fd_sc_hd__clkbuf_2 _12140_ (.A(_05932_),
    .X(_05949_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(_01367_),
    .A1(_04576_),
    .S(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__clkbuf_1 _12142_ (.A(_05950_),
    .X(_00024_));
 sky130_fd_sc_hd__nor2_1 _12143_ (.A(\core.mem_do_prefetch ),
    .B(\core.mem_do_rinst ),
    .Y(_05951_));
 sky130_fd_sc_hd__clkbuf_2 _12144_ (.A(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__clkbuf_2 _12145_ (.A(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__clkbuf_2 _12146_ (.A(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__inv_2 _12147_ (.A(\core.reg_out[17] ),
    .Y(_05955_));
 sky130_fd_sc_hd__nand2_2 _12148_ (.A(\core.latched_store ),
    .B(\core.latched_branch ),
    .Y(_05956_));
 sky130_fd_sc_hd__clkbuf_2 _12149_ (.A(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12150_ (.A(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_2 _12151_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__inv_2 _12152_ (.A(_05951_),
    .Y(_05960_));
 sky130_fd_sc_hd__clkbuf_2 _12153_ (.A(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__clkbuf_2 _12154_ (.A(_05956_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_2 _12155_ (.A(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__nand2_1 _12156_ (.A(_05963_),
    .B(\core.reg_next_pc[17] ),
    .Y(_05964_));
 sky130_fd_sc_hd__o211a_1 _12157_ (.A1(_05955_),
    .A2(_05959_),
    .B1(_05961_),
    .C1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__a21oi_1 _12158_ (.A1(_04904_),
    .A2(_05954_),
    .B1(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__nor2_1 _12159_ (.A(\core.mem_do_rdata ),
    .B(_05960_),
    .Y(_05967_));
 sky130_fd_sc_hd__inv_2 _12160_ (.A(_04371_),
    .Y(_05968_));
 sky130_fd_sc_hd__a211o_1 _12161_ (.A1(_05967_),
    .A2(_04370_),
    .B1(_04512_),
    .C1(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__inv_2 _12162_ (.A(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__inv_2 _12163_ (.A(net103),
    .Y(_05971_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_05970_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__clkbuf_2 _12165_ (.A(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__mux2_1 _12166_ (.A0(_05966_),
    .A1(net42),
    .S(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _12167_ (.A(_05974_),
    .X(_00037_));
 sky130_fd_sc_hd__inv_2 _12168_ (.A(\core.reg_out[18] ),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2_2 _12169_ (.A(_05962_),
    .B(\core.reg_next_pc[18] ),
    .Y(_05976_));
 sky130_fd_sc_hd__o211a_1 _12170_ (.A1(_05975_),
    .A2(_05959_),
    .B1(_05961_),
    .C1(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__a21oi_1 _12171_ (.A1(_04909_),
    .A2(_05954_),
    .B1(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__clkbuf_2 _12172_ (.A(_05972_),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(_05978_),
    .A1(net43),
    .S(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__buf_1 _12174_ (.A(_05980_),
    .X(_00038_));
 sky130_fd_sc_hd__inv_2 _12175_ (.A(\core.reg_out[19] ),
    .Y(_05981_));
 sky130_fd_sc_hd__clkbuf_4 _12176_ (.A(_05960_),
    .X(_05982_));
 sky130_fd_sc_hd__clkbuf_2 _12177_ (.A(_05956_),
    .X(_05983_));
 sky130_fd_sc_hd__nand2_1 _12178_ (.A(_05983_),
    .B(\core.reg_next_pc[19] ),
    .Y(_05984_));
 sky130_fd_sc_hd__o211a_1 _12179_ (.A1(_05981_),
    .A2(_05959_),
    .B1(_05982_),
    .C1(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__a21oi_2 _12180_ (.A1(_04911_),
    .A2(_05954_),
    .B1(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(_05986_),
    .A1(net44),
    .S(_05979_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_05987_),
    .X(_00039_));
 sky130_fd_sc_hd__inv_2 _12183_ (.A(\core.reg_out[20] ),
    .Y(_05988_));
 sky130_fd_sc_hd__clkbuf_2 _12184_ (.A(_05958_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_2 _12185_ (.A(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__nand2_1 _12186_ (.A(_05963_),
    .B(\core.reg_next_pc[20] ),
    .Y(_05991_));
 sky130_fd_sc_hd__o211a_1 _12187_ (.A1(_05988_),
    .A2(_05990_),
    .B1(_05982_),
    .C1(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__a21oi_1 _12188_ (.A1(_04917_),
    .A2(_05954_),
    .B1(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__mux2_1 _12189_ (.A0(_05993_),
    .A1(net45),
    .S(_05979_),
    .X(_05994_));
 sky130_fd_sc_hd__clkbuf_1 _12190_ (.A(_05994_),
    .X(_00040_));
 sky130_fd_sc_hd__inv_2 _12191_ (.A(\core.reg_out[21] ),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(_05957_),
    .B(\core.reg_next_pc[21] ),
    .Y(_05996_));
 sky130_fd_sc_hd__o211a_1 _12193_ (.A1(_05995_),
    .A2(_05990_),
    .B1(_05982_),
    .C1(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a21oi_1 _12194_ (.A1(_04916_),
    .A2(_05954_),
    .B1(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(_05998_),
    .A1(net46),
    .S(_05979_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _12196_ (.A(_05999_),
    .X(_00041_));
 sky130_fd_sc_hd__inv_2 _12197_ (.A(\core.reg_out[22] ),
    .Y(_06000_));
 sky130_fd_sc_hd__buf_6 _12198_ (.A(_05983_),
    .X(_06001_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(_06001_),
    .B(\core.reg_next_pc[22] ),
    .Y(_06002_));
 sky130_fd_sc_hd__o211a_1 _12200_ (.A1(_06000_),
    .A2(_05990_),
    .B1(_05982_),
    .C1(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__a21oi_1 _12201_ (.A1(_04924_),
    .A2(_05954_),
    .B1(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__mux2_1 _12202_ (.A0(_06004_),
    .A1(net47),
    .S(_05979_),
    .X(_06005_));
 sky130_fd_sc_hd__buf_1 _12203_ (.A(_06005_),
    .X(_00042_));
 sky130_fd_sc_hd__clkinv_4 _12204_ (.A(_05956_),
    .Y(_06006_));
 sky130_fd_sc_hd__buf_6 _12205_ (.A(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__buf_6 _12206_ (.A(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__buf_6 _12207_ (.A(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_2 _12208_ (.A(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_2 _12209_ (.A(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__nand2_2 _12210_ (.A(_05963_),
    .B(\core.reg_next_pc[23] ),
    .Y(_06012_));
 sky130_fd_sc_hd__a21bo_1 _12211_ (.A1(\core.reg_out[23] ),
    .A2(_06011_),
    .B1_N(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__mux2_1 _12212_ (.A0(_06013_),
    .A1(_04879_),
    .S(_05953_),
    .X(_06014_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(_06014_),
    .A1(net48),
    .S(_05979_),
    .X(_06015_));
 sky130_fd_sc_hd__clkbuf_1 _12214_ (.A(_06015_),
    .X(_00043_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05963_),
    .B(\core.reg_next_pc[24] ),
    .Y(_06016_));
 sky130_fd_sc_hd__a21bo_1 _12216_ (.A1(\core.reg_out[24] ),
    .A2(_06011_),
    .B1_N(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(_06017_),
    .A1(_04829_),
    .S(_05953_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_4 _12218_ (.A(_05972_),
    .X(_06019_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(_06018_),
    .A1(net49),
    .S(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _12220_ (.A(_06020_),
    .X(_00044_));
 sky130_fd_sc_hd__clkbuf_2 _12221_ (.A(_05960_),
    .X(_06021_));
 sky130_fd_sc_hd__nand2_1 _12222_ (.A(_06001_),
    .B(\core.reg_next_pc[25] ),
    .Y(_06022_));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__a21o_1 _12224_ (.A1(_06011_),
    .A2(\core.reg_out[25] ),
    .B1(_05952_),
    .X(_06024_));
 sky130_fd_sc_hd__o22a_1 _12225_ (.A1(\core.pcpi_rs1[25] ),
    .A2(_06021_),
    .B1(_06023_),
    .B2(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_06025_),
    .A1(net50),
    .S(_06019_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _12227_ (.A(_06026_),
    .X(_00045_));
 sky130_fd_sc_hd__nand2_1 _12228_ (.A(_06001_),
    .B(\core.reg_next_pc[26] ),
    .Y(_06027_));
 sky130_fd_sc_hd__inv_2 _12229_ (.A(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a21o_1 _12230_ (.A1(_06011_),
    .A2(\core.reg_out[26] ),
    .B1(_05952_),
    .X(_06029_));
 sky130_fd_sc_hd__o22a_1 _12231_ (.A1(\core.pcpi_rs1[26] ),
    .A2(_06021_),
    .B1(_06028_),
    .B2(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(_06030_),
    .A1(net51),
    .S(_06019_),
    .X(_06031_));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(_06031_),
    .X(_00046_));
 sky130_fd_sc_hd__clkbuf_2 _12234_ (.A(\core.pcpi_rs1[27] ),
    .X(_06032_));
 sky130_fd_sc_hd__nand2_2 _12235_ (.A(_05962_),
    .B(\core.reg_next_pc[27] ),
    .Y(_06033_));
 sky130_fd_sc_hd__inv_2 _12236_ (.A(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__inv_2 _12237_ (.A(\core.reg_out[27] ),
    .Y(_06035_));
 sky130_fd_sc_hd__o21ai_1 _12238_ (.A1(_06035_),
    .A2(_05959_),
    .B1(_05961_),
    .Y(_06036_));
 sky130_fd_sc_hd__o22a_1 _12239_ (.A1(_06032_),
    .A2(_06021_),
    .B1(_06034_),
    .B2(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(_06037_),
    .A1(net52),
    .S(_06019_),
    .X(_06038_));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(_06038_),
    .X(_00047_));
 sky130_fd_sc_hd__nand2_2 _12242_ (.A(_05957_),
    .B(\core.reg_next_pc[28] ),
    .Y(_06039_));
 sky130_fd_sc_hd__inv_2 _12243_ (.A(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__inv_2 _12244_ (.A(\core.reg_out[28] ),
    .Y(_06041_));
 sky130_fd_sc_hd__o21ai_2 _12245_ (.A1(_06041_),
    .A2(_05959_),
    .B1(_05961_),
    .Y(_06042_));
 sky130_fd_sc_hd__o22a_1 _12246_ (.A1(_04849_),
    .A2(_06021_),
    .B1(_06040_),
    .B2(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__mux2_1 _12247_ (.A0(_06043_),
    .A1(net53),
    .S(_06019_),
    .X(_06044_));
 sky130_fd_sc_hd__buf_1 _12248_ (.A(_06044_),
    .X(_00048_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_05958_),
    .B(\core.reg_next_pc[29] ),
    .Y(_06045_));
 sky130_fd_sc_hd__inv_2 _12250_ (.A(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__a21o_1 _12251_ (.A1(_06011_),
    .A2(\core.reg_out[29] ),
    .B1(_05952_),
    .X(_06047_));
 sky130_fd_sc_hd__o22a_1 _12252_ (.A1(_04856_),
    .A2(_06021_),
    .B1(_06046_),
    .B2(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(_06048_),
    .A1(net54),
    .S(_06019_),
    .X(_06049_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_06049_),
    .X(_00049_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(_05958_),
    .B(\core.reg_next_pc[30] ),
    .Y(_06050_));
 sky130_fd_sc_hd__inv_2 _12256_ (.A(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__inv_2 _12257_ (.A(\core.reg_out[30] ),
    .Y(_06052_));
 sky130_fd_sc_hd__o21ai_1 _12258_ (.A1(_06052_),
    .A2(_05959_),
    .B1(_05961_),
    .Y(_06053_));
 sky130_fd_sc_hd__o22a_1 _12259_ (.A1(_04845_),
    .A2(_05961_),
    .B1(_06051_),
    .B2(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__buf_4 _12260_ (.A(_05972_),
    .X(_06055_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(_06054_),
    .A1(net56),
    .S(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_06056_),
    .X(_00050_));
 sky130_fd_sc_hd__nand2_1 _12263_ (.A(_05958_),
    .B(\core.reg_next_pc[31] ),
    .Y(_06057_));
 sky130_fd_sc_hd__a21bo_1 _12264_ (.A1(\core.reg_out[31] ),
    .A2(_06011_),
    .B1_N(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__buf_4 _12265_ (.A(_05951_),
    .X(_06059_));
 sky130_fd_sc_hd__mux2_1 _12266_ (.A0(_06058_),
    .A1(\core.pcpi_rs1[31] ),
    .S(_06059_),
    .X(_06060_));
 sky130_fd_sc_hd__mux2_2 _12267_ (.A0(_06060_),
    .A1(net57),
    .S(_06055_),
    .X(_06061_));
 sky130_fd_sc_hd__buf_1 _12268_ (.A(_06061_),
    .X(_00051_));
 sky130_fd_sc_hd__nor2_2 _12269_ (.A(_04728_),
    .B(\core.decoded_imm[5] ),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_1 _12270_ (.A(_04728_),
    .B(\core.decoded_imm[5] ),
    .Y(_06063_));
 sky130_fd_sc_hd__inv_2 _12271_ (.A(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__nor2_1 _12272_ (.A(_06062_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_2 _12273_ (.A(_04723_),
    .B(\core.decoded_imm[4] ),
    .Y(_06066_));
 sky130_fd_sc_hd__or2_1 _12274_ (.A(_04723_),
    .B(\core.decoded_imm[4] ),
    .X(_06067_));
 sky130_fd_sc_hd__and3_1 _12275_ (.A(_06065_),
    .B(_06066_),
    .C(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(_04734_),
    .B(\core.decoded_imm[7] ),
    .Y(_06069_));
 sky130_fd_sc_hd__nand2_1 _12277_ (.A(_04734_),
    .B(\core.decoded_imm[7] ),
    .Y(_06070_));
 sky130_fd_sc_hd__and2b_1 _12278_ (.A_N(_06069_),
    .B(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__nor2_2 _12279_ (.A(_04737_),
    .B(\core.decoded_imm[6] ),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_1 _12280_ (.A(_04737_),
    .B(\core.decoded_imm[6] ),
    .Y(_06073_));
 sky130_fd_sc_hd__and2b_1 _12281_ (.A_N(_06072_),
    .B(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__and2_1 _12282_ (.A(_06071_),
    .B(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__nand2_1 _12283_ (.A(_06068_),
    .B(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand2_1 _12284_ (.A(\core.pcpi_rs1[0] ),
    .B(\core.decoded_imm[0] ),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_1 _12285_ (.A(_04688_),
    .B(_05021_),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_1 _12286_ (.A(\core.pcpi_rs1[1] ),
    .B(\core.decoded_imm[1] ),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2_1 _12287_ (.A(_06078_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__nor2_1 _12288_ (.A(_06077_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__inv_2 _12289_ (.A(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_1 _12290_ (.A(_06082_),
    .B(_06079_),
    .Y(_06083_));
 sky130_fd_sc_hd__or2_1 _12291_ (.A(\core.pcpi_rs1[3] ),
    .B(\core.decoded_imm[3] ),
    .X(_06084_));
 sky130_fd_sc_hd__nand2_1 _12292_ (.A(_04677_),
    .B(\core.decoded_imm[3] ),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_06084_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__inv_2 _12294_ (.A(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_1 _12295_ (.A(_04683_),
    .B(_05054_),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2_2 _12296_ (.A(\core.pcpi_rs1[2] ),
    .B(\core.decoded_imm[2] ),
    .Y(_06089_));
 sky130_fd_sc_hd__and2_1 _12297_ (.A(_06088_),
    .B(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__nand3_1 _12298_ (.A(_06083_),
    .B(_06087_),
    .C(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__o21a_1 _12299_ (.A1(_06089_),
    .A2(_06086_),
    .B1(_06085_),
    .X(_06092_));
 sky130_fd_sc_hd__nand2_1 _12300_ (.A(_06091_),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__inv_2 _12301_ (.A(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__o21a_1 _12302_ (.A1(_06066_),
    .A2(_06062_),
    .B1(_06063_),
    .X(_06095_));
 sky130_fd_sc_hd__inv_2 _12303_ (.A(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21ai_1 _12304_ (.A1(_06073_),
    .A2(_06069_),
    .B1(_06070_),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_2 _12305_ (.A1(_06075_),
    .A2(_06096_),
    .B1(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__o21ai_2 _12306_ (.A1(_06076_),
    .A2(_06094_),
    .B1(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nor2_1 _12307_ (.A(\core.pcpi_rs1[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_2 _12308_ (.A(\core.pcpi_rs1[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_06101_));
 sky130_fd_sc_hd__and2b_1 _12309_ (.A_N(_06100_),
    .B(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__nor2_1 _12310_ (.A(\core.pcpi_rs1[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_06103_));
 sky130_fd_sc_hd__nand2_1 _12311_ (.A(\core.pcpi_rs1[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_06104_));
 sky130_fd_sc_hd__nor2b_1 _12312_ (.A(_06103_),
    .B_N(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand2_1 _12313_ (.A(_06102_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__inv_2 _12314_ (.A(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__nor2_1 _12315_ (.A(\core.pcpi_rs1[15] ),
    .B(\core.decoded_imm[15] ),
    .Y(_06108_));
 sky130_fd_sc_hd__nand2_1 _12316_ (.A(\core.pcpi_rs1[15] ),
    .B(\core.decoded_imm[15] ),
    .Y(_06109_));
 sky130_fd_sc_hd__inv_2 _12317_ (.A(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__nor2_1 _12318_ (.A(_06108_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__inv_2 _12319_ (.A(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_1 _12320_ (.A(\core.pcpi_rs1[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_1 _12321_ (.A(\core.pcpi_rs1[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_06114_));
 sky130_fd_sc_hd__inv_2 _12322_ (.A(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__nor2_1 _12323_ (.A(_06113_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__inv_2 _12324_ (.A(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _12325_ (.A(_06112_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_1 _12326_ (.A(_06107_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__inv_2 _12327_ (.A(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__nor2_1 _12328_ (.A(\core.pcpi_rs1[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_06121_));
 sky130_fd_sc_hd__nand2_2 _12329_ (.A(\core.pcpi_rs1[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_06122_));
 sky130_fd_sc_hd__inv_2 _12330_ (.A(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__nor2_2 _12331_ (.A(_06121_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__nor2_1 _12332_ (.A(\core.pcpi_rs1[11] ),
    .B(\core.decoded_imm[11] ),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_8 _12333_ (.A(\core.pcpi_rs1[11] ),
    .B(\core.decoded_imm[11] ),
    .Y(_06126_));
 sky130_fd_sc_hd__inv_2 _12334_ (.A(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__nor2_2 _12335_ (.A(_06125_),
    .B(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_8 _12336_ (.A(_06124_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__inv_2 _12337_ (.A(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__inv_2 _12338_ (.A(\core.decoded_imm[8] ),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_1 _12339_ (.A(_04783_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(\core.pcpi_rs1[8] ),
    .B(\core.decoded_imm[8] ),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2_2 _12341_ (.A(_06132_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__nor2_1 _12342_ (.A(_04752_),
    .B(\core.decoded_imm[9] ),
    .Y(_06135_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(_04752_),
    .B(\core.decoded_imm[9] ),
    .Y(_06136_));
 sky130_fd_sc_hd__or2b_2 _12344_ (.A(_06135_),
    .B_N(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__nor2_2 _12345_ (.A(_06134_),
    .B(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__and3_1 _12346_ (.A(_06120_),
    .B(_06130_),
    .C(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_1 _12347_ (.A(_06099_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__inv_2 _12348_ (.A(_06128_),
    .Y(_06141_));
 sky130_fd_sc_hd__o21a_2 _12349_ (.A1(_06133_),
    .A2(_06135_),
    .B1(_06136_),
    .X(_06142_));
 sky130_fd_sc_hd__o221ai_4 _12350_ (.A1(_06122_),
    .A2(_06141_),
    .B1(_06129_),
    .B2(_06142_),
    .C1(_06126_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21a_1 _12351_ (.A1(_06101_),
    .A2(_06103_),
    .B1(_06104_),
    .X(_06144_));
 sky130_fd_sc_hd__o21a_1 _12352_ (.A1(_06114_),
    .A2(_06108_),
    .B1(_06109_),
    .X(_06145_));
 sky130_fd_sc_hd__o31ai_1 _12353_ (.A1(_06112_),
    .A2(_06117_),
    .A3(_06144_),
    .B1(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__a21oi_1 _12354_ (.A1(_06143_),
    .A2(_06120_),
    .B1(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__nand2_1 _12355_ (.A(_06140_),
    .B(_06147_),
    .Y(_06148_));
 sky130_fd_sc_hd__nor2_1 _12356_ (.A(_04879_),
    .B(\core.decoded_imm[23] ),
    .Y(_06149_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(_04879_),
    .B(\core.decoded_imm[23] ),
    .Y(_06150_));
 sky130_fd_sc_hd__and2b_1 _12358_ (.A_N(_06149_),
    .B(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__nor2_1 _12359_ (.A(\core.pcpi_rs1[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(\core.pcpi_rs1[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_06153_));
 sky130_fd_sc_hd__and2b_2 _12361_ (.A_N(_06152_),
    .B(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _12362_ (.A(_06151_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__nor2_1 _12363_ (.A(\core.pcpi_rs1[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_06156_));
 sky130_fd_sc_hd__nand2_1 _12364_ (.A(\core.pcpi_rs1[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_06157_));
 sky130_fd_sc_hd__inv_2 _12365_ (.A(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__or2_1 _12366_ (.A(_06156_),
    .B(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__inv_2 _12367_ (.A(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_2 _12368_ (.A(\core.pcpi_rs1[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_4 _12369_ (.A(\core.pcpi_rs1[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_06162_));
 sky130_fd_sc_hd__and2b_2 _12370_ (.A_N(_06161_),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__and3b_1 _12371_ (.A_N(_06155_),
    .B(_06160_),
    .C(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_1 _12372_ (.A(\core.pcpi_rs1[18] ),
    .B(\core.decoded_imm[18] ),
    .Y(_06165_));
 sky130_fd_sc_hd__nand2_1 _12373_ (.A(\core.pcpi_rs1[18] ),
    .B(\core.decoded_imm[18] ),
    .Y(_06166_));
 sky130_fd_sc_hd__and2b_1 _12374_ (.A_N(_06165_),
    .B(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__nor2_1 _12375_ (.A(\core.pcpi_rs1[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_06168_));
 sky130_fd_sc_hd__nand2_1 _12376_ (.A(\core.pcpi_rs1[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_06169_));
 sky130_fd_sc_hd__inv_2 _12377_ (.A(_06169_),
    .Y(_06170_));
 sky130_fd_sc_hd__nor2_2 _12378_ (.A(_06168_),
    .B(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_1 _12379_ (.A(_06167_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__nor2_1 _12380_ (.A(\core.pcpi_rs1[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _12381_ (.A(\core.pcpi_rs1[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_06174_));
 sky130_fd_sc_hd__and2b_1 _12382_ (.A_N(_06173_),
    .B(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__nor2_4 _12383_ (.A(\core.pcpi_rs1[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_06176_));
 sky130_fd_sc_hd__nand2_1 _12384_ (.A(\core.pcpi_rs1[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_06177_));
 sky130_fd_sc_hd__and2b_1 _12385_ (.A_N(_06176_),
    .B(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__nand2_1 _12386_ (.A(_06175_),
    .B(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__nor2_1 _12387_ (.A(_06172_),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__and2_4 _12388_ (.A(_06164_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__nand2_1 _12389_ (.A(_06148_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__inv_2 _12390_ (.A(_06171_),
    .Y(_06183_));
 sky130_fd_sc_hd__o21a_1 _12391_ (.A1(_06177_),
    .A2(_06173_),
    .B1(_06174_),
    .X(_06184_));
 sky130_fd_sc_hd__o221ai_4 _12392_ (.A1(_06183_),
    .A2(_06166_),
    .B1(_06184_),
    .B2(_06172_),
    .C1(_06169_),
    .Y(_06185_));
 sky130_fd_sc_hd__o21a_1 _12393_ (.A1(_06162_),
    .A2(_06156_),
    .B1(_06157_),
    .X(_06186_));
 sky130_fd_sc_hd__o221a_1 _12394_ (.A1(_06149_),
    .A2(_06153_),
    .B1(_06186_),
    .B2(_06155_),
    .C1(_06150_),
    .X(_06187_));
 sky130_fd_sc_hd__a21boi_1 _12395_ (.A1(_06164_),
    .A2(_06185_),
    .B1_N(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_2 _12396_ (.A(_06182_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__inv_2 _12397_ (.A(\core.decoded_imm[26] ),
    .Y(_06190_));
 sky130_fd_sc_hd__nand2_8 _12398_ (.A(_04819_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand2_1 _12399_ (.A(\core.pcpi_rs1[26] ),
    .B(\core.decoded_imm[26] ),
    .Y(_06192_));
 sky130_fd_sc_hd__and2_1 _12400_ (.A(_06191_),
    .B(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__nor2_1 _12401_ (.A(_06032_),
    .B(\core.decoded_imm[27] ),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_2 _12402_ (.A(_06032_),
    .B(\core.decoded_imm[27] ),
    .Y(_06195_));
 sky130_fd_sc_hd__and2b_1 _12403_ (.A_N(_06194_),
    .B(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__nor2_1 _12404_ (.A(\core.pcpi_rs1[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_8 _12405_ (.A(\core.pcpi_rs1[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_06198_));
 sky130_fd_sc_hd__and2b_1 _12406_ (.A_N(_06197_),
    .B(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__nor2_8 _12407_ (.A(_04829_),
    .B(\core.decoded_imm[24] ),
    .Y(_06200_));
 sky130_fd_sc_hd__nand2_1 _12408_ (.A(_04829_),
    .B(\core.decoded_imm[24] ),
    .Y(_06201_));
 sky130_fd_sc_hd__and2b_2 _12409_ (.A_N(_06200_),
    .B(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__and4_1 _12410_ (.A(_06193_),
    .B(_06196_),
    .C(_06199_),
    .D(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__nand2_1 _12411_ (.A(_06189_),
    .B(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__o21a_1 _12412_ (.A1(_06201_),
    .A2(_06197_),
    .B1(_06198_),
    .X(_06205_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_06196_),
    .B(_06193_),
    .Y(_06206_));
 sky130_fd_sc_hd__o221a_1 _12414_ (.A1(_06194_),
    .A2(_06192_),
    .B1(_06205_),
    .B2(_06206_),
    .C1(_06195_),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_1 _12415_ (.A(_06204_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nor2_2 _12416_ (.A(_04856_),
    .B(\core.decoded_imm[29] ),
    .Y(_06209_));
 sky130_fd_sc_hd__nand2_2 _12417_ (.A(_04856_),
    .B(\core.decoded_imm[29] ),
    .Y(_06210_));
 sky130_fd_sc_hd__and2b_2 _12418_ (.A_N(_06209_),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__nor2_1 _12419_ (.A(_04849_),
    .B(\core.decoded_imm[28] ),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_2 _12420_ (.A(_04849_),
    .B(\core.decoded_imm[28] ),
    .Y(_06213_));
 sky130_fd_sc_hd__and2b_1 _12421_ (.A_N(_06212_),
    .B(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__nand3_1 _12422_ (.A(_06208_),
    .B(_06211_),
    .C(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__o21a_1 _12423_ (.A1(_06213_),
    .A2(_06209_),
    .B1(_06210_),
    .X(_06216_));
 sky130_fd_sc_hd__nand2_2 _12424_ (.A(_06215_),
    .B(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__nand2_1 _12425_ (.A(_04843_),
    .B(_05519_),
    .Y(_06218_));
 sky130_fd_sc_hd__nand2_1 _12426_ (.A(_04845_),
    .B(\core.decoded_imm[30] ),
    .Y(_06219_));
 sky130_fd_sc_hd__and2_1 _12427_ (.A(_06218_),
    .B(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__nand2_1 _12428_ (.A(_06217_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__nand2_1 _12429_ (.A(_06221_),
    .B(_06219_),
    .Y(_06222_));
 sky130_fd_sc_hd__xor2_4 _12430_ (.A(\core.pcpi_rs1[31] ),
    .B(\core.decoded_imm[31] ),
    .X(_06223_));
 sky130_fd_sc_hd__nand2_1 _12431_ (.A(_06222_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__buf_4 _12432_ (.A(_04397_),
    .X(_06225_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12433_ (.A(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__inv_2 _12434_ (.A(_06223_),
    .Y(_06227_));
 sky130_fd_sc_hd__nand3_1 _12435_ (.A(_06221_),
    .B(_06219_),
    .C(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__nand3_1 _12436_ (.A(_06224_),
    .B(_06226_),
    .C(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__clkbuf_4 _12437_ (.A(_04506_),
    .X(_06230_));
 sky130_fd_sc_hd__nor2_2 _12438_ (.A(\core.instr_sra ),
    .B(\core.instr_srai ),
    .Y(_06231_));
 sky130_fd_sc_hd__nor2_1 _12439_ (.A(\core.instr_srl ),
    .B(\core.instr_srli ),
    .Y(_06232_));
 sky130_fd_sc_hd__nand2_1 _12440_ (.A(_06231_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__clkbuf_4 _12441_ (.A(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12442_ (.A(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(_06032_),
    .A1(_04845_),
    .S(_04481_),
    .X(_06236_));
 sky130_fd_sc_hd__or3b_1 _12444_ (.A(_06230_),
    .B(_06235_),
    .C_N(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__buf_2 _12445_ (.A(_00005_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_4 _12446_ (.A(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_2 _12447_ (.A(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__mux2_2 _12448_ (.A0(\core.cpuregs[12][31] ),
    .A1(\core.cpuregs[13][31] ),
    .S(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12449_ (.A(_06238_),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_2 _12450_ (.A(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\core.cpuregs[14][31] ),
    .A1(\core.cpuregs[15][31] ),
    .S(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__buf_2 _12452_ (.A(_00006_),
    .X(_06245_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12453_ (.A(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_2 _12454_ (.A(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(_06241_),
    .A1(_06244_),
    .S(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__mux2_1 _12456_ (.A0(\core.cpuregs[8][31] ),
    .A1(\core.cpuregs[9][31] ),
    .S(_06243_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_2 _12457_ (.A(_06242_),
    .X(_06250_));
 sky130_fd_sc_hd__mux2_1 _12458_ (.A0(\core.cpuregs[10][31] ),
    .A1(\core.cpuregs[11][31] ),
    .S(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(_06249_),
    .A1(_06251_),
    .S(_06247_),
    .X(_06252_));
 sky130_fd_sc_hd__inv_2 _12460_ (.A(_00007_),
    .Y(_06253_));
 sky130_fd_sc_hd__clkbuf_2 _12461_ (.A(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(_06248_),
    .A1(_06252_),
    .S(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_2 _12463_ (.A(_06242_),
    .X(_06256_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(\core.cpuregs[24][31] ),
    .A1(\core.cpuregs[25][31] ),
    .S(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\core.cpuregs[26][31] ),
    .A1(\core.cpuregs[27][31] ),
    .S(_06250_),
    .X(_06258_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(_06257_),
    .A1(_06258_),
    .S(_06247_),
    .X(_06259_));
 sky130_fd_sc_hd__buf_4 _12467_ (.A(_06242_),
    .X(_06260_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(\core.cpuregs[28][31] ),
    .A1(\core.cpuregs[29][31] ),
    .S(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__clkbuf_4 _12469_ (.A(_06242_),
    .X(_06262_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\core.cpuregs[30][31] ),
    .A1(\core.cpuregs[31][31] ),
    .S(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_4 _12471_ (.A(_06246_),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(_06261_),
    .A1(_06263_),
    .S(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__buf_2 _12473_ (.A(_00007_),
    .X(_06266_));
 sky130_fd_sc_hd__mux2_8 _12474_ (.A0(_06259_),
    .A1(_06265_),
    .S(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__buf_4 _12475_ (.A(_00009_),
    .X(_06268_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(_06255_),
    .A1(_06267_),
    .S(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__mux2_1 _12477_ (.A0(\core.cpuregs[0][31] ),
    .A1(\core.cpuregs[1][31] ),
    .S(_06260_),
    .X(_06270_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(\core.cpuregs[2][31] ),
    .A1(\core.cpuregs[3][31] ),
    .S(_06262_),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(_06270_),
    .A1(_06271_),
    .S(_06264_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_2 _12480_ (.A(_06242_),
    .X(_06273_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(\core.cpuregs[6][31] ),
    .A1(\core.cpuregs[7][31] ),
    .S(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_4 _12482_ (.A(_06238_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_2 _12483_ (.A(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(\core.cpuregs[4][31] ),
    .A1(\core.cpuregs[5][31] ),
    .S(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__inv_2 _12485_ (.A(_00006_),
    .Y(_06278_));
 sky130_fd_sc_hd__clkbuf_2 _12486_ (.A(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(_06274_),
    .A1(_06277_),
    .S(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(_06272_),
    .A1(_06280_),
    .S(_06266_),
    .X(_06281_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(\core.cpuregs[16][31] ),
    .A1(\core.cpuregs[17][31] ),
    .S(_06273_),
    .X(_06282_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(\core.cpuregs[18][31] ),
    .A1(\core.cpuregs[19][31] ),
    .S(_06276_),
    .X(_06283_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(_06282_),
    .A1(_06283_),
    .S(_06264_),
    .X(_06284_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(\core.cpuregs[22][31] ),
    .A1(\core.cpuregs[23][31] ),
    .S(_06262_),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(\core.cpuregs[20][31] ),
    .A1(\core.cpuregs[21][31] ),
    .S(_06276_),
    .X(_06286_));
 sky130_fd_sc_hd__mux2_1 _12494_ (.A0(_06285_),
    .A1(_06286_),
    .S(_06279_),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_2 _12495_ (.A(_00007_),
    .X(_06288_));
 sky130_fd_sc_hd__mux2_4 _12496_ (.A0(_06284_),
    .A1(_06287_),
    .S(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(_06281_),
    .A1(_06289_),
    .S(_06268_),
    .X(_06290_));
 sky130_fd_sc_hd__inv_2 _12498_ (.A(_00008_),
    .Y(_06291_));
 sky130_fd_sc_hd__clkbuf_4 _12499_ (.A(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__buf_2 _12500_ (.A(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(_06269_),
    .A1(_06290_),
    .S(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__nor3_1 _12502_ (.A(\core.decoded_imm_j[17] ),
    .B(\core.decoded_imm_j[18] ),
    .C(\core.decoded_imm_j[19] ),
    .Y(_06295_));
 sky130_fd_sc_hd__inv_2 _12503_ (.A(\core.decoded_imm_j[15] ),
    .Y(_06296_));
 sky130_fd_sc_hd__inv_2 _12504_ (.A(\core.decoded_imm_j[16] ),
    .Y(_06297_));
 sky130_fd_sc_hd__a31o_1 _12505_ (.A1(_06295_),
    .A2(_06296_),
    .A3(_06297_),
    .B1(\core.is_lui_auipc_jal ),
    .X(_06298_));
 sky130_fd_sc_hd__inv_2 _12506_ (.A(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_06294_),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__buf_1 _12508_ (.A(\core.instr_lui ),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_4 _12509_ (.A(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__inv_2 _12510_ (.A(\core.reg_pc[31] ),
    .Y(_06303_));
 sky130_fd_sc_hd__inv_2 _12511_ (.A(\core.is_lui_auipc_jal ),
    .Y(_06304_));
 sky130_fd_sc_hd__buf_1 _12512_ (.A(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__or3_1 _12513_ (.A(_06302_),
    .B(_06303_),
    .C(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__nand2_1 _12514_ (.A(_06300_),
    .B(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__nor2_1 _12515_ (.A(\core.cpu_state[4] ),
    .B(_04397_),
    .Y(_06308_));
 sky130_fd_sc_hd__buf_4 _12516_ (.A(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__nand2_1 _12517_ (.A(_06307_),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand3_2 _12518_ (.A(_06229_),
    .B(_06237_),
    .C(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__inv_2 _12519_ (.A(_04389_),
    .Y(_06312_));
 sky130_fd_sc_hd__or4_1 _12520_ (.A(\core.instr_sll ),
    .B(\core.instr_slli ),
    .C(_06233_),
    .D(_04484_),
    .X(_06313_));
 sky130_fd_sc_hd__nor2_1 _12521_ (.A(\core.cpu_state[2] ),
    .B(\core.cpu_state[4] ),
    .Y(_06314_));
 sky130_fd_sc_hd__inv_2 _12522_ (.A(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__nor2_2 _12523_ (.A(_04396_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nor2_8 _12524_ (.A(_04512_),
    .B(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__and3_1 _12525_ (.A(_06313_),
    .B(_04590_),
    .C(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__nand2_2 _12526_ (.A(_06318_),
    .B(_04398_),
    .Y(_06319_));
 sky130_fd_sc_hd__inv_2 _12527_ (.A(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__and3_1 _12528_ (.A(_04400_),
    .B(_06312_),
    .C(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__o21a_2 _12529_ (.A1(_04484_),
    .A2(_06231_),
    .B1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__nand2_8 _12530_ (.A(_06311_),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__or2_1 _12531_ (.A(_04838_),
    .B(_06322_),
    .X(_06324_));
 sky130_fd_sc_hd__nand2_1 _12532_ (.A(_06323_),
    .B(_06324_),
    .Y(_00052_));
 sky130_fd_sc_hd__buf_1 _12533_ (.A(_04513_),
    .X(_06325_));
 sky130_fd_sc_hd__buf_1 _12534_ (.A(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12535_ (.A(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__nor2_1 _12536_ (.A(\core.count_cycle[0] ),
    .B(_06327_),
    .Y(_00053_));
 sky130_fd_sc_hd__or2_1 _12537_ (.A(\core.count_cycle[0] ),
    .B(\core.count_cycle[1] ),
    .X(_06328_));
 sky130_fd_sc_hd__clkbuf_2 _12538_ (.A(_04451_),
    .X(_06329_));
 sky130_fd_sc_hd__nand2_1 _12539_ (.A(\core.count_cycle[0] ),
    .B(\core.count_cycle[1] ),
    .Y(_06330_));
 sky130_fd_sc_hd__and3_1 _12540_ (.A(_06328_),
    .B(_06329_),
    .C(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__buf_1 _12541_ (.A(_06331_),
    .X(_00054_));
 sky130_fd_sc_hd__inv_2 _12542_ (.A(_06330_),
    .Y(_06332_));
 sky130_fd_sc_hd__or2_1 _12543_ (.A(\core.count_cycle[2] ),
    .B(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__nand2_1 _12544_ (.A(_06332_),
    .B(\core.count_cycle[2] ),
    .Y(_06334_));
 sky130_fd_sc_hd__and3_1 _12545_ (.A(_06333_),
    .B(_06329_),
    .C(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__buf_1 _12546_ (.A(_06335_),
    .X(_00055_));
 sky130_fd_sc_hd__inv_2 _12547_ (.A(\core.count_cycle[3] ),
    .Y(_06336_));
 sky130_fd_sc_hd__nor2_1 _12548_ (.A(_06336_),
    .B(_06334_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _12549_ (.A(_06334_),
    .B(_06336_),
    .Y(_06338_));
 sky130_fd_sc_hd__and3b_1 _12550_ (.A_N(_06337_),
    .B(_04451_),
    .C(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__buf_1 _12551_ (.A(_06339_),
    .X(_00056_));
 sky130_fd_sc_hd__or2_1 _12552_ (.A(\core.count_cycle[4] ),
    .B(_06337_),
    .X(_06340_));
 sky130_fd_sc_hd__nand2_1 _12553_ (.A(_06337_),
    .B(\core.count_cycle[4] ),
    .Y(_06341_));
 sky130_fd_sc_hd__and3_1 _12554_ (.A(_06340_),
    .B(_06329_),
    .C(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__buf_1 _12555_ (.A(_06342_),
    .X(_00057_));
 sky130_fd_sc_hd__inv_2 _12556_ (.A(_06341_),
    .Y(_06343_));
 sky130_fd_sc_hd__nor2_1 _12557_ (.A(\core.count_cycle[5] ),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_06343_),
    .B(\core.count_cycle[5] ),
    .Y(_06345_));
 sky130_fd_sc_hd__or3b_2 _12559_ (.A(_06325_),
    .B(_06344_),
    .C_N(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__inv_2 _12560_ (.A(_06346_),
    .Y(_00058_));
 sky130_fd_sc_hd__inv_2 _12561_ (.A(\core.count_cycle[6] ),
    .Y(_06347_));
 sky130_fd_sc_hd__or2_2 _12562_ (.A(_06347_),
    .B(_06345_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(_06345_),
    .B(_06347_),
    .Y(_06349_));
 sky130_fd_sc_hd__and3_1 _12564_ (.A(_06348_),
    .B(_06329_),
    .C(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__buf_1 _12565_ (.A(_06350_),
    .X(_00059_));
 sky130_fd_sc_hd__inv_2 _12566_ (.A(\core.count_cycle[7] ),
    .Y(_06351_));
 sky130_fd_sc_hd__or2_2 _12567_ (.A(_06351_),
    .B(_06348_),
    .X(_06352_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(_06348_),
    .B(_06351_),
    .Y(_06353_));
 sky130_fd_sc_hd__and3_1 _12569_ (.A(_06352_),
    .B(_06329_),
    .C(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _12570_ (.A(_06354_),
    .X(_00060_));
 sky130_fd_sc_hd__inv_2 _12571_ (.A(\core.count_cycle[8] ),
    .Y(_06355_));
 sky130_fd_sc_hd__or2_2 _12572_ (.A(_06355_),
    .B(_06352_),
    .X(_06356_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12573_ (.A(_04388_),
    .X(_06357_));
 sky130_fd_sc_hd__clkbuf_2 _12574_ (.A(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__nand2_1 _12575_ (.A(_06352_),
    .B(_06355_),
    .Y(_06359_));
 sky130_fd_sc_hd__and3_1 _12576_ (.A(_06356_),
    .B(_06358_),
    .C(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__buf_1 _12577_ (.A(_06360_),
    .X(_00061_));
 sky130_fd_sc_hd__inv_2 _12578_ (.A(\core.count_cycle[9] ),
    .Y(_06361_));
 sky130_fd_sc_hd__nor2_2 _12579_ (.A(_06361_),
    .B(_06356_),
    .Y(_06362_));
 sky130_fd_sc_hd__inv_2 _12580_ (.A(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand2_1 _12581_ (.A(_06356_),
    .B(_06361_),
    .Y(_06364_));
 sky130_fd_sc_hd__and3_1 _12582_ (.A(_06363_),
    .B(_06358_),
    .C(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _12583_ (.A(_06365_),
    .X(_00062_));
 sky130_fd_sc_hd__inv_2 _12584_ (.A(\core.count_cycle[10] ),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_1 _12585_ (.A(_06363_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__nand2_4 _12586_ (.A(_06362_),
    .B(\core.count_cycle[10] ),
    .Y(_06368_));
 sky130_fd_sc_hd__and3_1 _12587_ (.A(_06367_),
    .B(_06358_),
    .C(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__buf_1 _12588_ (.A(_06369_),
    .X(_00063_));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(\core.count_cycle[11] ),
    .B(_06368_),
    .X(_06370_));
 sky130_fd_sc_hd__nand2_1 _12590_ (.A(_06368_),
    .B(\core.count_cycle[11] ),
    .Y(_06371_));
 sky130_fd_sc_hd__clkbuf_2 _12591_ (.A(_06326_),
    .X(_06372_));
 sky130_fd_sc_hd__a21oi_1 _12592_ (.A1(_06370_),
    .A2(_06371_),
    .B1(_06372_),
    .Y(_00064_));
 sky130_fd_sc_hd__and4_1 _12593_ (.A(_06362_),
    .B(\core.count_cycle[10] ),
    .C(\core.count_cycle[11] ),
    .D(\core.count_cycle[12] ),
    .X(_06373_));
 sky130_fd_sc_hd__inv_2 _12594_ (.A(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__a31o_1 _12595_ (.A1(_06362_),
    .A2(\core.count_cycle[10] ),
    .A3(\core.count_cycle[11] ),
    .B1(\core.count_cycle[12] ),
    .X(_06375_));
 sky130_fd_sc_hd__and3_1 _12596_ (.A(_06374_),
    .B(_06358_),
    .C(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__buf_1 _12597_ (.A(_06376_),
    .X(_00065_));
 sky130_fd_sc_hd__or2_1 _12598_ (.A(\core.count_cycle[13] ),
    .B(_06373_),
    .X(_06377_));
 sky130_fd_sc_hd__nand2_1 _12599_ (.A(_06373_),
    .B(\core.count_cycle[13] ),
    .Y(_06378_));
 sky130_fd_sc_hd__and3_1 _12600_ (.A(_06377_),
    .B(_06358_),
    .C(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_06379_),
    .X(_00066_));
 sky130_fd_sc_hd__inv_2 _12602_ (.A(\core.count_cycle[14] ),
    .Y(_06380_));
 sky130_fd_sc_hd__nor2_1 _12603_ (.A(_06380_),
    .B(_06378_),
    .Y(_06381_));
 sky130_fd_sc_hd__or2_1 _12604_ (.A(_06325_),
    .B(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__a21oi_1 _12605_ (.A1(_06380_),
    .A2(_06378_),
    .B1(_06382_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _12606_ (.A(\core.count_cycle[15] ),
    .Y(_06383_));
 sky130_fd_sc_hd__or2_1 _12607_ (.A(_06383_),
    .B(_06381_),
    .X(_06384_));
 sky130_fd_sc_hd__nand2_1 _12608_ (.A(_06381_),
    .B(_06383_),
    .Y(_06385_));
 sky130_fd_sc_hd__clkbuf_2 _12609_ (.A(_06326_),
    .X(_06386_));
 sky130_fd_sc_hd__a21oi_1 _12610_ (.A1(_06384_),
    .A2(_06385_),
    .B1(_06386_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_2 _12611_ (.A(\core.count_cycle[12] ),
    .B(\core.count_cycle[13] ),
    .Y(_06387_));
 sky130_fd_sc_hd__or4b_1 _12612_ (.A(_06355_),
    .B(_06361_),
    .C(_06366_),
    .D_N(\core.count_cycle[11] ),
    .X(_06388_));
 sky130_fd_sc_hd__or4_1 _12613_ (.A(_06380_),
    .B(_06383_),
    .C(_06387_),
    .D(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nor2_1 _12614_ (.A(_06352_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__clkbuf_2 _12615_ (.A(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(\core.count_cycle[16] ),
    .B(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__nand2_1 _12617_ (.A(_06391_),
    .B(\core.count_cycle[16] ),
    .Y(_06393_));
 sky130_fd_sc_hd__and3_1 _12618_ (.A(_06392_),
    .B(_06358_),
    .C(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _12619_ (.A(_06394_),
    .X(_00069_));
 sky130_fd_sc_hd__or2_2 _12620_ (.A(\core.count_cycle[17] ),
    .B(_06393_),
    .X(_06395_));
 sky130_fd_sc_hd__nand2_1 _12621_ (.A(_06393_),
    .B(\core.count_cycle[17] ),
    .Y(_06396_));
 sky130_fd_sc_hd__a21oi_2 _12622_ (.A1(_06395_),
    .A2(_06396_),
    .B1(_06386_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _12623_ (.A(\core.count_cycle[16] ),
    .B(\core.count_cycle[17] ),
    .Y(_06397_));
 sky130_fd_sc_hd__inv_2 _12624_ (.A(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__and2_1 _12625_ (.A(_06391_),
    .B(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__or2_1 _12626_ (.A(\core.count_cycle[18] ),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_2 _12627_ (.A(_06357_),
    .X(_06401_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(_06399_),
    .B(\core.count_cycle[18] ),
    .Y(_06402_));
 sky130_fd_sc_hd__and3_1 _12629_ (.A(_06400_),
    .B(_06401_),
    .C(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__buf_1 _12630_ (.A(_06403_),
    .X(_00071_));
 sky130_fd_sc_hd__or2_1 _12631_ (.A(\core.count_cycle[19] ),
    .B(_06402_),
    .X(_06404_));
 sky130_fd_sc_hd__nand2_2 _12632_ (.A(_06402_),
    .B(\core.count_cycle[19] ),
    .Y(_06405_));
 sky130_fd_sc_hd__a21oi_1 _12633_ (.A1(_06404_),
    .A2(_06405_),
    .B1(_06386_),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_2 _12634_ (.A(\core.count_cycle[20] ),
    .Y(_06406_));
 sky130_fd_sc_hd__and3_1 _12635_ (.A(_06398_),
    .B(\core.count_cycle[18] ),
    .C(\core.count_cycle[19] ),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_1 _12636_ (.A(_06391_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__or2_1 _12637_ (.A(_06406_),
    .B(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__nand2_1 _12638_ (.A(_06408_),
    .B(_06406_),
    .Y(_06410_));
 sky130_fd_sc_hd__and3_1 _12639_ (.A(_06409_),
    .B(_06401_),
    .C(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _12640_ (.A(_06411_),
    .X(_00073_));
 sky130_fd_sc_hd__or2_1 _12641_ (.A(\core.count_cycle[21] ),
    .B(_06409_),
    .X(_06412_));
 sky130_fd_sc_hd__nand2_1 _12642_ (.A(_06409_),
    .B(\core.count_cycle[21] ),
    .Y(_06413_));
 sky130_fd_sc_hd__a21oi_1 _12643_ (.A1(_06412_),
    .A2(_06413_),
    .B1(_06386_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _12644_ (.A(\core.count_cycle[22] ),
    .Y(_06414_));
 sky130_fd_sc_hd__nand2_1 _12645_ (.A(\core.count_cycle[20] ),
    .B(\core.count_cycle[21] ),
    .Y(_06415_));
 sky130_fd_sc_hd__or2_1 _12646_ (.A(_06415_),
    .B(_06408_),
    .X(_06416_));
 sky130_fd_sc_hd__nor2_1 _12647_ (.A(_06414_),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__inv_2 _12648_ (.A(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(_06416_),
    .B(_06414_),
    .Y(_06419_));
 sky130_fd_sc_hd__and3_1 _12650_ (.A(_06418_),
    .B(_06401_),
    .C(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__buf_1 _12651_ (.A(_06420_),
    .X(_00075_));
 sky130_fd_sc_hd__or2_1 _12652_ (.A(\core.count_cycle[23] ),
    .B(_06418_),
    .X(_06421_));
 sky130_fd_sc_hd__nand2_1 _12653_ (.A(_06418_),
    .B(\core.count_cycle[23] ),
    .Y(_06422_));
 sky130_fd_sc_hd__a21oi_2 _12654_ (.A1(_06421_),
    .A2(_06422_),
    .B1(_06386_),
    .Y(_00076_));
 sky130_fd_sc_hd__and4b_1 _12655_ (.A_N(_06415_),
    .B(_06407_),
    .C(\core.count_cycle[22] ),
    .D(\core.count_cycle[23] ),
    .X(_06423_));
 sky130_fd_sc_hd__nand2_2 _12656_ (.A(_06390_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__inv_2 _12657_ (.A(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _12658_ (.A(_06425_),
    .B(\core.count_cycle[24] ),
    .Y(_06426_));
 sky130_fd_sc_hd__inv_2 _12659_ (.A(\core.count_cycle[24] ),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(_06424_),
    .B(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__and3_1 _12661_ (.A(_06426_),
    .B(_06401_),
    .C(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__clkbuf_1 _12662_ (.A(_06429_),
    .X(_00077_));
 sky130_fd_sc_hd__or2_1 _12663_ (.A(\core.count_cycle[25] ),
    .B(_06426_),
    .X(_06430_));
 sky130_fd_sc_hd__nand2_1 _12664_ (.A(_06426_),
    .B(\core.count_cycle[25] ),
    .Y(_06431_));
 sky130_fd_sc_hd__a21oi_1 _12665_ (.A1(_06430_),
    .A2(_06431_),
    .B1(_06386_),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_2 _12666_ (.A(\core.count_cycle[26] ),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_1 _12667_ (.A(\core.count_cycle[24] ),
    .B(\core.count_cycle[25] ),
    .Y(_06433_));
 sky130_fd_sc_hd__or3_2 _12668_ (.A(_06432_),
    .B(_06433_),
    .C(_06424_),
    .X(_06434_));
 sky130_fd_sc_hd__o21ai_1 _12669_ (.A1(_06433_),
    .A2(_06424_),
    .B1(_06432_),
    .Y(_06435_));
 sky130_fd_sc_hd__and3_1 _12670_ (.A(_06434_),
    .B(_06401_),
    .C(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_06436_),
    .X(_00079_));
 sky130_fd_sc_hd__or2_2 _12672_ (.A(\core.count_cycle[27] ),
    .B(_06434_),
    .X(_06437_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(_06434_),
    .B(\core.count_cycle[27] ),
    .Y(_06438_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12674_ (.A(_06326_),
    .X(_06439_));
 sky130_fd_sc_hd__a21oi_1 _12675_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06439_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _12676_ (.A(\core.count_cycle[28] ),
    .Y(_06440_));
 sky130_fd_sc_hd__and4_1 _12677_ (.A(\core.count_cycle[24] ),
    .B(\core.count_cycle[25] ),
    .C(\core.count_cycle[26] ),
    .D(\core.count_cycle[27] ),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_1 _12678_ (.A(_06425_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__or2_1 _12679_ (.A(_06440_),
    .B(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__nand2_1 _12680_ (.A(_06442_),
    .B(_06440_),
    .Y(_06444_));
 sky130_fd_sc_hd__and3_1 _12681_ (.A(_06443_),
    .B(_06401_),
    .C(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _12682_ (.A(_06445_),
    .X(_00081_));
 sky130_fd_sc_hd__or2_1 _12683_ (.A(\core.count_cycle[29] ),
    .B(_06443_),
    .X(_06446_));
 sky130_fd_sc_hd__nand2_1 _12684_ (.A(_06443_),
    .B(\core.count_cycle[29] ),
    .Y(_06447_));
 sky130_fd_sc_hd__a21oi_1 _12685_ (.A1(_06446_),
    .A2(_06447_),
    .B1(_06439_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(\core.count_cycle[28] ),
    .B(\core.count_cycle[29] ),
    .Y(_06448_));
 sky130_fd_sc_hd__nor2_1 _12687_ (.A(_06448_),
    .B(_06442_),
    .Y(_06449_));
 sky130_fd_sc_hd__or2_1 _12688_ (.A(\core.count_cycle[30] ),
    .B(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_2 _12689_ (.A(_06357_),
    .X(_06451_));
 sky130_fd_sc_hd__nand2_1 _12690_ (.A(_06449_),
    .B(\core.count_cycle[30] ),
    .Y(_06452_));
 sky130_fd_sc_hd__and3_1 _12691_ (.A(_06450_),
    .B(_06451_),
    .C(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__buf_1 _12692_ (.A(_06453_),
    .X(_00083_));
 sky130_fd_sc_hd__or2_1 _12693_ (.A(\core.count_cycle[31] ),
    .B(_06452_),
    .X(_06454_));
 sky130_fd_sc_hd__nand2_1 _12694_ (.A(_06452_),
    .B(\core.count_cycle[31] ),
    .Y(_06455_));
 sky130_fd_sc_hd__a21oi_1 _12695_ (.A1(_06454_),
    .A2(_06455_),
    .B1(_06439_),
    .Y(_00084_));
 sky130_fd_sc_hd__and4_1 _12696_ (.A(\core.count_cycle[28] ),
    .B(\core.count_cycle[29] ),
    .C(\core.count_cycle[30] ),
    .D(\core.count_cycle[31] ),
    .X(_06456_));
 sky130_fd_sc_hd__and3_1 _12697_ (.A(_06425_),
    .B(_06441_),
    .C(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__or2_1 _12698_ (.A(\core.count_cycle[32] ),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__nand2_1 _12699_ (.A(_06457_),
    .B(\core.count_cycle[32] ),
    .Y(_06459_));
 sky130_fd_sc_hd__and3_1 _12700_ (.A(_06458_),
    .B(_06451_),
    .C(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _12701_ (.A(_06460_),
    .X(_00085_));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(\core.count_cycle[33] ),
    .B(_06459_),
    .X(_06461_));
 sky130_fd_sc_hd__nand2_1 _12703_ (.A(_06459_),
    .B(\core.count_cycle[33] ),
    .Y(_06462_));
 sky130_fd_sc_hd__a21oi_1 _12704_ (.A1(_06461_),
    .A2(_06462_),
    .B1(_06439_),
    .Y(_00086_));
 sky130_fd_sc_hd__and3_1 _12705_ (.A(_06423_),
    .B(_06441_),
    .C(_06456_),
    .X(_06463_));
 sky130_fd_sc_hd__nand2_1 _12706_ (.A(_06391_),
    .B(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__inv_2 _12707_ (.A(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand2_1 _12708_ (.A(\core.count_cycle[32] ),
    .B(\core.count_cycle[33] ),
    .Y(_06466_));
 sky130_fd_sc_hd__inv_2 _12709_ (.A(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__nand2_2 _12710_ (.A(_06465_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__nor2_1 _12711_ (.A(_05040_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__or2_1 _12712_ (.A(_06325_),
    .B(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__a21oi_1 _12713_ (.A1(_05040_),
    .A2(_06468_),
    .B1(_06470_),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _12714_ (.A(\core.count_cycle[35] ),
    .Y(_06471_));
 sky130_fd_sc_hd__or2_1 _12715_ (.A(_06471_),
    .B(_06469_),
    .X(_06472_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(_06469_),
    .B(_06471_),
    .Y(_06473_));
 sky130_fd_sc_hd__a21oi_1 _12717_ (.A1(_06472_),
    .A2(_06473_),
    .B1(_06439_),
    .Y(_00088_));
 sky130_fd_sc_hd__and3_1 _12718_ (.A(_06467_),
    .B(\core.count_cycle[34] ),
    .C(\core.count_cycle[35] ),
    .X(_06474_));
 sky130_fd_sc_hd__nand2_1 _12719_ (.A(_06465_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__inv_2 _12720_ (.A(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__or2_1 _12721_ (.A(\core.count_cycle[36] ),
    .B(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__nand2_1 _12722_ (.A(_06476_),
    .B(\core.count_cycle[36] ),
    .Y(_06478_));
 sky130_fd_sc_hd__and3_1 _12723_ (.A(_06477_),
    .B(_06451_),
    .C(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__buf_1 _12724_ (.A(_06479_),
    .X(_00089_));
 sky130_fd_sc_hd__or2_1 _12725_ (.A(\core.count_cycle[37] ),
    .B(_06478_),
    .X(_06480_));
 sky130_fd_sc_hd__nand2_1 _12726_ (.A(_06478_),
    .B(\core.count_cycle[37] ),
    .Y(_06481_));
 sky130_fd_sc_hd__a21oi_1 _12727_ (.A1(_06480_),
    .A2(_06481_),
    .B1(_06439_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_1 _12728_ (.A(\core.count_cycle[36] ),
    .B(\core.count_cycle[37] ),
    .Y(_06482_));
 sky130_fd_sc_hd__nor2_1 _12729_ (.A(_06482_),
    .B(_06475_),
    .Y(_06483_));
 sky130_fd_sc_hd__or2_1 _12730_ (.A(\core.count_cycle[38] ),
    .B(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__nand2_1 _12731_ (.A(_06483_),
    .B(\core.count_cycle[38] ),
    .Y(_06485_));
 sky130_fd_sc_hd__and3_1 _12732_ (.A(_06484_),
    .B(_06451_),
    .C(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__buf_1 _12733_ (.A(_06486_),
    .X(_00091_));
 sky130_fd_sc_hd__or2_1 _12734_ (.A(\core.count_cycle[39] ),
    .B(_06485_),
    .X(_06487_));
 sky130_fd_sc_hd__nand2_1 _12735_ (.A(_06485_),
    .B(\core.count_cycle[39] ),
    .Y(_06488_));
 sky130_fd_sc_hd__buf_2 _12736_ (.A(_06326_),
    .X(_06489_));
 sky130_fd_sc_hd__a21oi_1 _12737_ (.A1(_06487_),
    .A2(_06488_),
    .B1(_06489_),
    .Y(_00092_));
 sky130_fd_sc_hd__and4_1 _12738_ (.A(\core.count_cycle[36] ),
    .B(\core.count_cycle[37] ),
    .C(\core.count_cycle[38] ),
    .D(\core.count_cycle[39] ),
    .X(_06490_));
 sky130_fd_sc_hd__and2_1 _12739_ (.A(_06490_),
    .B(_06474_),
    .X(_06491_));
 sky130_fd_sc_hd__nand2_2 _12740_ (.A(_06465_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__or2_1 _12741_ (.A(\core.count_cycle[40] ),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__nand2_1 _12742_ (.A(_06492_),
    .B(\core.count_cycle[40] ),
    .Y(_06494_));
 sky130_fd_sc_hd__a21oi_1 _12743_ (.A1(_06493_),
    .A2(_06494_),
    .B1(_06489_),
    .Y(_00093_));
 sky130_fd_sc_hd__or3b_1 _12744_ (.A(\core.count_cycle[41] ),
    .B(_06492_),
    .C_N(\core.count_cycle[40] ),
    .X(_06495_));
 sky130_fd_sc_hd__inv_2 _12745_ (.A(\core.count_cycle[41] ),
    .Y(_06496_));
 sky130_fd_sc_hd__a31o_1 _12746_ (.A1(_06465_),
    .A2(\core.count_cycle[40] ),
    .A3(_06491_),
    .B1(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__a21oi_1 _12747_ (.A1(_06495_),
    .A2(_06497_),
    .B1(_06489_),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _12748_ (.A(\core.count_cycle[42] ),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_2 _12749_ (.A(\core.count_cycle[40] ),
    .B(\core.count_cycle[41] ),
    .Y(_06499_));
 sky130_fd_sc_hd__nor2_1 _12750_ (.A(_06499_),
    .B(_06492_),
    .Y(_06500_));
 sky130_fd_sc_hd__or2_1 _12751_ (.A(_06498_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(_06500_),
    .B(_06498_),
    .Y(_06502_));
 sky130_fd_sc_hd__a21oi_1 _12753_ (.A1(_06501_),
    .A2(_06502_),
    .B1(_06489_),
    .Y(_00095_));
 sky130_fd_sc_hd__inv_2 _12754_ (.A(\core.count_cycle[43] ),
    .Y(_06503_));
 sky130_fd_sc_hd__a21oi_1 _12755_ (.A1(_06500_),
    .A2(\core.count_cycle[42] ),
    .B1(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__and3_1 _12756_ (.A(_06500_),
    .B(\core.count_cycle[42] ),
    .C(_06503_),
    .X(_06505_));
 sky130_fd_sc_hd__buf_2 _12757_ (.A(_04451_),
    .X(_06506_));
 sky130_fd_sc_hd__o21a_1 _12758_ (.A1(_06504_),
    .A2(_06505_),
    .B1(_06506_),
    .X(_00096_));
 sky130_fd_sc_hd__inv_2 _12759_ (.A(\core.count_cycle[44] ),
    .Y(_06507_));
 sky130_fd_sc_hd__or3_1 _12760_ (.A(_06498_),
    .B(_06503_),
    .C(_06499_),
    .X(_06508_));
 sky130_fd_sc_hd__nor2_2 _12761_ (.A(_06508_),
    .B(_06492_),
    .Y(_06509_));
 sky130_fd_sc_hd__or2_1 _12762_ (.A(_06507_),
    .B(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__nand2_1 _12763_ (.A(_06509_),
    .B(_06507_),
    .Y(_06511_));
 sky130_fd_sc_hd__a21oi_1 _12764_ (.A1(_06510_),
    .A2(_06511_),
    .B1(_06489_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _12765_ (.A(_06509_),
    .B(\core.count_cycle[44] ),
    .Y(_06512_));
 sky130_fd_sc_hd__or2_1 _12766_ (.A(\core.count_cycle[45] ),
    .B(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__nand2_1 _12767_ (.A(_06512_),
    .B(\core.count_cycle[45] ),
    .Y(_06514_));
 sky130_fd_sc_hd__a21oi_1 _12768_ (.A1(_06513_),
    .A2(_06514_),
    .B1(_06489_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _12769_ (.A(\core.count_cycle[44] ),
    .B(\core.count_cycle[45] ),
    .Y(_06515_));
 sky130_fd_sc_hd__inv_2 _12770_ (.A(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_1 _12771_ (.A(_06509_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__or2_1 _12772_ (.A(\core.count_cycle[46] ),
    .B(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__nand2_1 _12773_ (.A(_06517_),
    .B(\core.count_cycle[46] ),
    .Y(_06519_));
 sky130_fd_sc_hd__buf_1 _12774_ (.A(_06325_),
    .X(_06520_));
 sky130_fd_sc_hd__buf_2 _12775_ (.A(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__a21oi_1 _12776_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06521_),
    .Y(_00099_));
 sky130_fd_sc_hd__and2_1 _12777_ (.A(_06509_),
    .B(_06516_),
    .X(_06522_));
 sky130_fd_sc_hd__nand3b_2 _12778_ (.A_N(\core.count_cycle[47] ),
    .B(_06522_),
    .C(\core.count_cycle[46] ),
    .Y(_06523_));
 sky130_fd_sc_hd__inv_2 _12779_ (.A(\core.count_cycle[46] ),
    .Y(_06524_));
 sky130_fd_sc_hd__o21ai_1 _12780_ (.A1(_06524_),
    .A2(_06517_),
    .B1(\core.count_cycle[47] ),
    .Y(_06525_));
 sky130_fd_sc_hd__a21oi_1 _12781_ (.A1(_06523_),
    .A2(_06525_),
    .B1(_06521_),
    .Y(_00100_));
 sky130_fd_sc_hd__and3_1 _12782_ (.A(_06516_),
    .B(\core.count_cycle[46] ),
    .C(\core.count_cycle[47] ),
    .X(_06526_));
 sky130_fd_sc_hd__and3b_1 _12783_ (.A_N(_06508_),
    .B(_06491_),
    .C(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__and3_1 _12784_ (.A(_06390_),
    .B(_06463_),
    .C(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__clkbuf_2 _12785_ (.A(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__inv_2 _12786_ (.A(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__or2_1 _12787_ (.A(\core.count_cycle[48] ),
    .B(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__nand2_1 _12788_ (.A(_06530_),
    .B(\core.count_cycle[48] ),
    .Y(_06532_));
 sky130_fd_sc_hd__a21oi_1 _12789_ (.A1(_06531_),
    .A2(_06532_),
    .B1(_06521_),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _12790_ (.A(\core.count_cycle[49] ),
    .Y(_06533_));
 sky130_fd_sc_hd__a21oi_1 _12791_ (.A1(_06529_),
    .A2(\core.count_cycle[48] ),
    .B1(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__and3_1 _12792_ (.A(_06529_),
    .B(\core.count_cycle[48] ),
    .C(_06533_),
    .X(_06535_));
 sky130_fd_sc_hd__o21a_1 _12793_ (.A1(_06534_),
    .A2(_06535_),
    .B1(_06506_),
    .X(_00102_));
 sky130_fd_sc_hd__inv_2 _12794_ (.A(\core.count_cycle[50] ),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _12795_ (.A(\core.count_cycle[48] ),
    .B(\core.count_cycle[49] ),
    .Y(_06537_));
 sky130_fd_sc_hd__nor2_1 _12796_ (.A(_06537_),
    .B(_06530_),
    .Y(_06538_));
 sky130_fd_sc_hd__or2_1 _12797_ (.A(_06536_),
    .B(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__nand2_1 _12798_ (.A(_06538_),
    .B(_06536_),
    .Y(_06540_));
 sky130_fd_sc_hd__a21oi_1 _12799_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06521_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _12800_ (.A(_06538_),
    .B(\core.count_cycle[50] ),
    .Y(_06541_));
 sky130_fd_sc_hd__or2_1 _12801_ (.A(\core.count_cycle[51] ),
    .B(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_06541_),
    .B(\core.count_cycle[51] ),
    .Y(_06543_));
 sky130_fd_sc_hd__a21oi_1 _12803_ (.A1(_06542_),
    .A2(_06543_),
    .B1(_06521_),
    .Y(_00104_));
 sky130_fd_sc_hd__or3b_1 _12804_ (.A(_06536_),
    .B(_06537_),
    .C_N(\core.count_cycle[51] ),
    .X(_06544_));
 sky130_fd_sc_hd__inv_2 _12805_ (.A(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_2 _12806_ (.A(_06529_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__or2_1 _12807_ (.A(\core.count_cycle[52] ),
    .B(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(_06546_),
    .B(\core.count_cycle[52] ),
    .Y(_06548_));
 sky130_fd_sc_hd__a21oi_1 _12809_ (.A1(_06547_),
    .A2(_06548_),
    .B1(_06521_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand3_1 _12810_ (.A(_06529_),
    .B(\core.count_cycle[52] ),
    .C(_06545_),
    .Y(_06549_));
 sky130_fd_sc_hd__or2_1 _12811_ (.A(\core.count_cycle[53] ),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__nand2_1 _12812_ (.A(_06549_),
    .B(\core.count_cycle[53] ),
    .Y(_06551_));
 sky130_fd_sc_hd__clkbuf_2 _12813_ (.A(_06520_),
    .X(_06552_));
 sky130_fd_sc_hd__a21oi_1 _12814_ (.A1(_06550_),
    .A2(_06551_),
    .B1(_06552_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_2 _12815_ (.A(\core.count_cycle[52] ),
    .B(\core.count_cycle[53] ),
    .Y(_06553_));
 sky130_fd_sc_hd__nor2_1 _12816_ (.A(_06553_),
    .B(_06546_),
    .Y(_06554_));
 sky130_fd_sc_hd__or2_1 _12817_ (.A(\core.count_cycle[54] ),
    .B(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nand2_1 _12818_ (.A(_06554_),
    .B(\core.count_cycle[54] ),
    .Y(_06556_));
 sky130_fd_sc_hd__and3_1 _12819_ (.A(_06555_),
    .B(_06451_),
    .C(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__clkbuf_1 _12820_ (.A(_06557_),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _12821_ (.A(_06556_),
    .B(\core.count_cycle[55] ),
    .Y(_06558_));
 sky130_fd_sc_hd__nand3b_1 _12822_ (.A_N(\core.count_cycle[55] ),
    .B(_06554_),
    .C(\core.count_cycle[54] ),
    .Y(_06559_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_06558_),
    .A2(_06559_),
    .B1(_06552_),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _12824_ (.A(\core.count_cycle[56] ),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_1 _12825_ (.A(\core.count_cycle[54] ),
    .B(\core.count_cycle[55] ),
    .Y(_06561_));
 sky130_fd_sc_hd__nor3_2 _12826_ (.A(_06553_),
    .B(_06561_),
    .C(_06544_),
    .Y(_06562_));
 sky130_fd_sc_hd__and4_2 _12827_ (.A(_06391_),
    .B(_06463_),
    .C(_06527_),
    .D(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__or2_1 _12828_ (.A(_06560_),
    .B(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__nand2_1 _12829_ (.A(_06563_),
    .B(_06560_),
    .Y(_06565_));
 sky130_fd_sc_hd__a21oi_1 _12830_ (.A1(_06564_),
    .A2(_06565_),
    .B1(_06552_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand2_1 _12831_ (.A(_06563_),
    .B(\core.count_cycle[56] ),
    .Y(_06566_));
 sky130_fd_sc_hd__or2_1 _12832_ (.A(\core.count_cycle[57] ),
    .B(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(_06566_),
    .B(\core.count_cycle[57] ),
    .Y(_06568_));
 sky130_fd_sc_hd__a21oi_1 _12834_ (.A1(_06567_),
    .A2(_06568_),
    .B1(_06552_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _12835_ (.A(\core.count_cycle[56] ),
    .B(\core.count_cycle[57] ),
    .Y(_06569_));
 sky130_fd_sc_hd__inv_2 _12836_ (.A(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__nand2_1 _12837_ (.A(_06563_),
    .B(_06570_),
    .Y(_06571_));
 sky130_fd_sc_hd__inv_2 _12838_ (.A(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__inv_2 _12839_ (.A(\core.count_cycle[58] ),
    .Y(_06573_));
 sky130_fd_sc_hd__nand2_1 _12840_ (.A(_06572_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_1 _12841_ (.A(_06571_),
    .B(\core.count_cycle[58] ),
    .Y(_06575_));
 sky130_fd_sc_hd__a21oi_1 _12842_ (.A1(_06574_),
    .A2(_06575_),
    .B1(_06552_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand3b_1 _12843_ (.A_N(\core.count_cycle[59] ),
    .B(_06572_),
    .C(\core.count_cycle[58] ),
    .Y(_06576_));
 sky130_fd_sc_hd__o21ai_2 _12844_ (.A1(_06573_),
    .A2(_06571_),
    .B1(\core.count_cycle[59] ),
    .Y(_06577_));
 sky130_fd_sc_hd__a21oi_1 _12845_ (.A1(_06576_),
    .A2(_06577_),
    .B1(_06552_),
    .Y(_00112_));
 sky130_fd_sc_hd__and3_1 _12846_ (.A(_06570_),
    .B(\core.count_cycle[58] ),
    .C(\core.count_cycle[59] ),
    .X(_06578_));
 sky130_fd_sc_hd__nand3_4 _12847_ (.A(_06529_),
    .B(_06562_),
    .C(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__or2_1 _12848_ (.A(\core.count_cycle[60] ),
    .B(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(_06579_),
    .B(\core.count_cycle[60] ),
    .Y(_06581_));
 sky130_fd_sc_hd__clkbuf_2 _12850_ (.A(_06520_),
    .X(_06582_));
 sky130_fd_sc_hd__a21oi_1 _12851_ (.A1(_06580_),
    .A2(_06581_),
    .B1(_06582_),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _12852_ (.A(\core.count_cycle[60] ),
    .Y(_06583_));
 sky130_fd_sc_hd__nor2_1 _12853_ (.A(_06583_),
    .B(_06579_),
    .Y(_06584_));
 sky130_fd_sc_hd__nand2b_1 _12854_ (.A_N(\core.count_cycle[61] ),
    .B(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__o21ai_1 _12855_ (.A1(_06583_),
    .A2(_06579_),
    .B1(\core.count_cycle[61] ),
    .Y(_06586_));
 sky130_fd_sc_hd__a21oi_1 _12856_ (.A1(_06585_),
    .A2(_06586_),
    .B1(_06582_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _12857_ (.A(\core.count_cycle[60] ),
    .B(\core.count_cycle[61] ),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2_1 _12858_ (.A(_06587_),
    .B(_06579_),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2b_1 _12859_ (.A_N(\core.count_cycle[62] ),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__o21ai_1 _12860_ (.A1(_06587_),
    .A2(_06579_),
    .B1(\core.count_cycle[62] ),
    .Y(_06590_));
 sky130_fd_sc_hd__a21oi_1 _12861_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06582_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _12862_ (.A(_06588_),
    .B(\core.count_cycle[62] ),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _12863_ (.A(_06591_),
    .B(\core.count_cycle[63] ),
    .Y(_06592_));
 sky130_fd_sc_hd__nand3b_1 _12864_ (.A_N(\core.count_cycle[63] ),
    .B(_06588_),
    .C(\core.count_cycle[62] ),
    .Y(_06593_));
 sky130_fd_sc_hd__a21oi_1 _12865_ (.A1(_06592_),
    .A2(_06593_),
    .B1(_06582_),
    .Y(_00116_));
 sky130_fd_sc_hd__clkbuf_2 _12866_ (.A(_06006_),
    .X(_06594_));
 sky130_fd_sc_hd__buf_2 _12867_ (.A(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__inv_2 _12868_ (.A(\core.latched_stalu ),
    .Y(_06596_));
 sky130_fd_sc_hd__clkbuf_2 _12869_ (.A(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__nand2_1 _12870_ (.A(_06597_),
    .B(\core.reg_out[1] ),
    .Y(_06598_));
 sky130_fd_sc_hd__buf_6 _12871_ (.A(\core.latched_stalu ),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_2 _12872_ (.A(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__clkbuf_2 _12873_ (.A(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nand2_1 _12874_ (.A(_06601_),
    .B(\core.alu_out_q[1] ),
    .Y(_06602_));
 sky130_fd_sc_hd__nand3_1 _12875_ (.A(_06595_),
    .B(_06598_),
    .C(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__or2b_2 _12876_ (.A(\core.reg_next_pc[1] ),
    .B_N(_05962_),
    .X(_06604_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(_06603_),
    .B(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__inv_2 _12878_ (.A(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__buf_1 _12879_ (.A(\core.instr_jal ),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_1 _12880_ (.A(\core.decoder_trigger ),
    .B(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__inv_2 _12881_ (.A(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__o21ai_1 _12882_ (.A1(_04578_),
    .A2(_06608_),
    .B1(_06605_),
    .Y(_06610_));
 sky130_fd_sc_hd__nand2_1 _12883_ (.A(_06610_),
    .B(_04391_),
    .Y(_06611_));
 sky130_fd_sc_hd__a31o_1 _12884_ (.A1(_05942_),
    .A2(_06606_),
    .A3(_06609_),
    .B1(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__nand2_1 _12885_ (.A(_04500_),
    .B(\core.reg_next_pc[1] ),
    .Y(_06613_));
 sky130_fd_sc_hd__a21oi_1 _12886_ (.A1(_06612_),
    .A2(_06613_),
    .B1(_06582_),
    .Y(_00117_));
 sky130_fd_sc_hd__nor2_1 _12887_ (.A(_04391_),
    .B(_04513_),
    .Y(_06614_));
 sky130_fd_sc_hd__buf_2 _12888_ (.A(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__buf_4 _12889_ (.A(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12890_ (.A(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__nand3_2 _12891_ (.A(_06603_),
    .B(_05942_),
    .C(_06604_),
    .Y(_06618_));
 sky130_fd_sc_hd__nand2_1 _12892_ (.A(_06596_),
    .B(\core.reg_out[2] ),
    .Y(_06619_));
 sky130_fd_sc_hd__buf_6 _12893_ (.A(\core.latched_stalu ),
    .X(_06620_));
 sky130_fd_sc_hd__nand2_1 _12894_ (.A(_06620_),
    .B(\core.alu_out_q[2] ),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(_06619_),
    .B(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_06622_),
    .B(_06006_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_1 _12897_ (.A(_05956_),
    .B(\core.reg_next_pc[2] ),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_1 _12898_ (.A(_06623_),
    .B(_06624_),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_1 _12899_ (.A(_06625_),
    .B(\core.decoded_imm_j[2] ),
    .Y(_06626_));
 sky130_fd_sc_hd__nand3_2 _12900_ (.A(_06623_),
    .B(_04579_),
    .C(_06624_),
    .Y(_06627_));
 sky130_fd_sc_hd__nand2_1 _12901_ (.A(_06626_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__or2_1 _12902_ (.A(_06618_),
    .B(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__nand2_1 _12903_ (.A(_06628_),
    .B(_06618_),
    .Y(_06630_));
 sky130_fd_sc_hd__buf_1 _12904_ (.A(\core.decoder_trigger ),
    .X(_06631_));
 sky130_fd_sc_hd__buf_1 _12905_ (.A(\core.instr_jal ),
    .X(_06632_));
 sky130_fd_sc_hd__o21ai_1 _12906_ (.A1(_06632_),
    .A2(_06625_),
    .B1(_06631_),
    .Y(_06633_));
 sky130_fd_sc_hd__o21a_1 _12907_ (.A1(_06631_),
    .A2(_06625_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__a31o_1 _12908_ (.A1(_06629_),
    .A2(_06609_),
    .A3(_06630_),
    .B1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__inv_2 _12909_ (.A(_04457_),
    .Y(_06636_));
 sky130_fd_sc_hd__clkbuf_4 _12910_ (.A(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__clkbuf_2 _12911_ (.A(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__a22o_1 _12912_ (.A1(\core.reg_next_pc[2] ),
    .A2(_06617_),
    .B1(_06635_),
    .B2(_06638_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _12913_ (.A(_06596_),
    .B(\core.reg_out[3] ),
    .Y(_06639_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(_06620_),
    .B(\core.alu_out_q[3] ),
    .Y(_06640_));
 sky130_fd_sc_hd__nand2_4 _12915_ (.A(_06639_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_1 _12916_ (.A(_06641_),
    .B(_06006_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand2_2 _12917_ (.A(_05956_),
    .B(\core.reg_next_pc[3] ),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_1 _12918_ (.A(_06642_),
    .B(_06643_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(_06644_),
    .B(_04575_),
    .Y(_06645_));
 sky130_fd_sc_hd__inv_2 _12920_ (.A(\core.decoded_imm_j[3] ),
    .Y(_06646_));
 sky130_fd_sc_hd__nand3_1 _12921_ (.A(_06642_),
    .B(_06646_),
    .C(_06643_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2_1 _12922_ (.A(_06645_),
    .B(_06647_),
    .Y(_06648_));
 sky130_fd_sc_hd__inv_2 _12923_ (.A(_06627_),
    .Y(_06649_));
 sky130_fd_sc_hd__o21ai_2 _12924_ (.A1(_06618_),
    .A2(_06649_),
    .B1(_06626_),
    .Y(_06650_));
 sky130_fd_sc_hd__inv_2 _12925_ (.A(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__or2_2 _12926_ (.A(_06648_),
    .B(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__nand2_1 _12927_ (.A(_06651_),
    .B(_06648_),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_1 _12928_ (.A(_06652_),
    .B(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_1 _12929_ (.A(_06625_),
    .B(_06644_),
    .Y(_06655_));
 sky130_fd_sc_hd__inv_2 _12930_ (.A(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__inv_2 _12931_ (.A(\core.instr_jal ),
    .Y(_06657_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12932_ (.A(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(_06654_),
    .A1(_06656_),
    .S(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12934_ (.A(_06631_),
    .X(_06660_));
 sky130_fd_sc_hd__nand2_1 _12935_ (.A(_06659_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__buf_2 _12936_ (.A(_06636_),
    .X(_06662_));
 sky130_fd_sc_hd__or2b_1 _12937_ (.A(_06644_),
    .B_N(_06633_),
    .X(_06663_));
 sky130_fd_sc_hd__clkbuf_2 _12938_ (.A(_06615_),
    .X(_06664_));
 sky130_fd_sc_hd__a32o_1 _12939_ (.A1(_06661_),
    .A2(_06662_),
    .A3(_06663_),
    .B1(net111),
    .B2(_06664_),
    .X(_00119_));
 sky130_fd_sc_hd__buf_2 _12940_ (.A(_06658_),
    .X(_06665_));
 sky130_fd_sc_hd__nand2_1 _12941_ (.A(_06597_),
    .B(\core.reg_out[4] ),
    .Y(_06666_));
 sky130_fd_sc_hd__buf_6 _12942_ (.A(_06620_),
    .X(_06667_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_06667_),
    .B(\core.alu_out_q[4] ),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_1 _12944_ (.A(_06666_),
    .B(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand2_1 _12945_ (.A(_06669_),
    .B(_06594_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_2 _12946_ (.A(_05962_),
    .B(\core.reg_next_pc[4] ),
    .Y(_06671_));
 sky130_fd_sc_hd__nand2_1 _12947_ (.A(_06670_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__or2_1 _12948_ (.A(_06672_),
    .B(_06656_),
    .X(_06673_));
 sky130_fd_sc_hd__nand2_1 _12949_ (.A(_06656_),
    .B(_06672_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand2_1 _12950_ (.A(_06672_),
    .B(_04576_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand3b_2 _12951_ (.A_N(\core.decoded_imm_j[4] ),
    .B(_06670_),
    .C(_06671_),
    .Y(_06676_));
 sky130_fd_sc_hd__nand2_1 _12952_ (.A(_06675_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__a31o_1 _12953_ (.A1(_06652_),
    .A2(_06645_),
    .A3(_06677_),
    .B1(_06657_),
    .X(_06678_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_06652_),
    .A2(_06645_),
    .B1(_06677_),
    .X(_06679_));
 sky130_fd_sc_hd__nor2b_1 _12955_ (.A(_06678_),
    .B_N(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__a31o_1 _12956_ (.A1(_06665_),
    .A2(_06673_),
    .A3(_06674_),
    .B1(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__clkbuf_2 _12957_ (.A(_04501_),
    .X(_06682_));
 sky130_fd_sc_hd__clkbuf_2 _12958_ (.A(_06682_),
    .X(_06683_));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(_06681_),
    .A1(_06672_),
    .S(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12960_ (.A(_06636_),
    .X(_06685_));
 sky130_fd_sc_hd__nand2_1 _12961_ (.A(_06664_),
    .B(\core.reg_next_pc[4] ),
    .Y(_06686_));
 sky130_fd_sc_hd__a21bo_1 _12962_ (.A1(_06684_),
    .A2(_06685_),
    .B1_N(_06686_),
    .X(_00120_));
 sky130_fd_sc_hd__nor2_1 _12963_ (.A(_06648_),
    .B(_06677_),
    .Y(_06687_));
 sky130_fd_sc_hd__nand2_1 _12964_ (.A(_06650_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__inv_2 _12965_ (.A(_06676_),
    .Y(_06689_));
 sky130_fd_sc_hd__o21a_1 _12966_ (.A1(_06645_),
    .A2(_06689_),
    .B1(_06675_),
    .X(_06690_));
 sky130_fd_sc_hd__nand2_1 _12967_ (.A(_06688_),
    .B(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__inv_2 _12968_ (.A(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_1 _12969_ (.A(_06597_),
    .B(\core.reg_out[5] ),
    .Y(_06693_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(_06599_),
    .B(\core.alu_out_q[5] ),
    .Y(_06694_));
 sky130_fd_sc_hd__nand2_1 _12971_ (.A(_06693_),
    .B(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_1 _12972_ (.A(_06695_),
    .B(_06007_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_1 _12973_ (.A(_05983_),
    .B(\core.reg_next_pc[5] ),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_4 _12974_ (.A(_06696_),
    .B(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__nand2_2 _12975_ (.A(_06698_),
    .B(\core.decoded_imm_j[5] ),
    .Y(_06699_));
 sky130_fd_sc_hd__nand3b_1 _12976_ (.A_N(\core.decoded_imm_j[5] ),
    .B(_06696_),
    .C(_06697_),
    .Y(_06700_));
 sky130_fd_sc_hd__nand2_2 _12977_ (.A(_06699_),
    .B(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand2_1 _12978_ (.A(_06692_),
    .B(_06701_),
    .Y(_06702_));
 sky130_fd_sc_hd__clkbuf_2 _12979_ (.A(_06607_),
    .X(_06703_));
 sky130_fd_sc_hd__inv_2 _12980_ (.A(_06701_),
    .Y(_06704_));
 sky130_fd_sc_hd__nand2_1 _12981_ (.A(_06691_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__inv_2 _12982_ (.A(_06698_),
    .Y(_06706_));
 sky130_fd_sc_hd__nor2_1 _12983_ (.A(_06706_),
    .B(_06674_),
    .Y(_06707_));
 sky130_fd_sc_hd__inv_2 _12984_ (.A(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand2_1 _12985_ (.A(_06674_),
    .B(_06706_),
    .Y(_06709_));
 sky130_fd_sc_hd__and3_1 _12986_ (.A(_06708_),
    .B(_06658_),
    .C(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a31o_1 _12987_ (.A1(_06702_),
    .A2(_06703_),
    .A3(_06705_),
    .B1(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__mux2_1 _12988_ (.A0(_06711_),
    .A1(_06698_),
    .S(_06683_),
    .X(_06712_));
 sky130_fd_sc_hd__a22o_1 _12989_ (.A1(\core.reg_next_pc[5] ),
    .A2(_06617_),
    .B1(_06712_),
    .B2(_06638_),
    .X(_00121_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(_06597_),
    .B(\core.reg_out[6] ),
    .Y(_06713_));
 sky130_fd_sc_hd__nand2_1 _12991_ (.A(_06599_),
    .B(\core.alu_out_q[6] ),
    .Y(_06714_));
 sky130_fd_sc_hd__nand2_2 _12992_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__nand2_2 _12993_ (.A(_06715_),
    .B(_06007_),
    .Y(_06716_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(_05983_),
    .B(\core.reg_next_pc[6] ),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_4 _12995_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__or2_1 _12996_ (.A(_06718_),
    .B(_06707_),
    .X(_06719_));
 sky130_fd_sc_hd__nand2_1 _12997_ (.A(_06707_),
    .B(_06718_),
    .Y(_06720_));
 sky130_fd_sc_hd__and2_1 _12998_ (.A(_06720_),
    .B(_06657_),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_1 _12999_ (.A(_06718_),
    .B(\core.decoded_imm_j[6] ),
    .Y(_06722_));
 sky130_fd_sc_hd__inv_2 _13000_ (.A(\core.decoded_imm_j[6] ),
    .Y(_06723_));
 sky130_fd_sc_hd__nand3_1 _13001_ (.A(_06716_),
    .B(_06723_),
    .C(_06717_),
    .Y(_06724_));
 sky130_fd_sc_hd__nand2_1 _13002_ (.A(_06722_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(_06725_),
    .Y(_06726_));
 sky130_fd_sc_hd__nand2_1 _13004_ (.A(_06705_),
    .B(_06699_),
    .Y(_06727_));
 sky130_fd_sc_hd__xor2_1 _13005_ (.A(_06726_),
    .B(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__a22o_1 _13006_ (.A1(_06719_),
    .A2(_06721_),
    .B1(_06728_),
    .B2(_06703_),
    .X(_06729_));
 sky130_fd_sc_hd__mux2_1 _13007_ (.A0(_06729_),
    .A1(_06718_),
    .S(_06683_),
    .X(_06730_));
 sky130_fd_sc_hd__a22o_1 _13008_ (.A1(net122),
    .A2(_06617_),
    .B1(_06730_),
    .B2(_06638_),
    .X(_00122_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13009_ (.A(_06632_),
    .X(_06731_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(_06597_),
    .B(\core.reg_out[7] ),
    .Y(_06732_));
 sky130_fd_sc_hd__nand2_1 _13011_ (.A(_06599_),
    .B(\core.alu_out_q[7] ),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_2 _13012_ (.A(_06732_),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand2_2 _13013_ (.A(_06734_),
    .B(_06007_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_1 _13014_ (.A(_05983_),
    .B(\core.reg_next_pc[7] ),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_2 _13015_ (.A(_06735_),
    .B(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_2 _13016_ (.A(_06718_),
    .B(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__nor2_1 _13017_ (.A(_06738_),
    .B(_06708_),
    .Y(_06739_));
 sky130_fd_sc_hd__and3_1 _13018_ (.A(_06720_),
    .B(_06736_),
    .C(_06735_),
    .X(_06740_));
 sky130_fd_sc_hd__nand2_1 _13019_ (.A(_06737_),
    .B(\core.decoded_imm_j[7] ),
    .Y(_06741_));
 sky130_fd_sc_hd__nand3b_1 _13020_ (.A_N(\core.decoded_imm_j[7] ),
    .B(_06735_),
    .C(_06736_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _13021_ (.A(_06741_),
    .B(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__inv_2 _13022_ (.A(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__nand2_1 _13023_ (.A(_06704_),
    .B(_06726_),
    .Y(_06745_));
 sky130_fd_sc_hd__inv_2 _13024_ (.A(_06724_),
    .Y(_06746_));
 sky130_fd_sc_hd__o21ai_1 _13025_ (.A1(_06699_),
    .A2(_06746_),
    .B1(_06722_),
    .Y(_06747_));
 sky130_fd_sc_hd__o21bai_1 _13026_ (.A1(_06745_),
    .A2(_06692_),
    .B1_N(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__or2_1 _13027_ (.A(_06744_),
    .B(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__nand2_1 _13028_ (.A(_06748_),
    .B(_06744_),
    .Y(_06750_));
 sky130_fd_sc_hd__nand3_1 _13029_ (.A(_06749_),
    .B(_06731_),
    .C(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__o31ai_1 _13030_ (.A1(_06731_),
    .A2(_06739_),
    .A3(_06740_),
    .B1(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(_06752_),
    .A1(_06737_),
    .S(_06683_),
    .X(_06753_));
 sky130_fd_sc_hd__a22o_1 _13032_ (.A1(\core.reg_next_pc[7] ),
    .A2(_06617_),
    .B1(_06753_),
    .B2(_06638_),
    .X(_00123_));
 sky130_fd_sc_hd__buf_6 _13033_ (.A(_06620_),
    .X(_06754_));
 sky130_fd_sc_hd__inv_2 _13034_ (.A(\core.reg_out[8] ),
    .Y(_06755_));
 sky130_fd_sc_hd__nand2_1 _13035_ (.A(_06754_),
    .B(\core.alu_out_q[8] ),
    .Y(_06756_));
 sky130_fd_sc_hd__o21ai_2 _13036_ (.A1(_06754_),
    .A2(_06755_),
    .B1(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(_06757_),
    .B(_06007_),
    .Y(_06758_));
 sky130_fd_sc_hd__nand2_1 _13038_ (.A(_05983_),
    .B(\core.reg_next_pc[8] ),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _13039_ (.A(_06758_),
    .B(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_1 _13040_ (.A(_06760_),
    .B(\core.decoded_imm_j[8] ),
    .Y(_06761_));
 sky130_fd_sc_hd__inv_2 _13041_ (.A(\core.decoded_imm_j[8] ),
    .Y(_06762_));
 sky130_fd_sc_hd__nand3_1 _13042_ (.A(_06758_),
    .B(_06762_),
    .C(_06759_),
    .Y(_06763_));
 sky130_fd_sc_hd__nand2_1 _13043_ (.A(_06761_),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__inv_2 _13044_ (.A(_06764_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_1 _13045_ (.A(_06750_),
    .B(_06741_),
    .Y(_06766_));
 sky130_fd_sc_hd__xor2_1 _13046_ (.A(_06765_),
    .B(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__nor2_1 _13047_ (.A(_06760_),
    .B(_06739_),
    .Y(_06768_));
 sky130_fd_sc_hd__inv_2 _13048_ (.A(_06738_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand3_2 _13049_ (.A(_06707_),
    .B(_06769_),
    .C(_06760_),
    .Y(_06770_));
 sky130_fd_sc_hd__and3b_1 _13050_ (.A_N(_06768_),
    .B(_06658_),
    .C(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a21o_1 _13051_ (.A1(_06767_),
    .A2(_06703_),
    .B1(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(_06772_),
    .A1(_06760_),
    .S(_06682_),
    .X(_06773_));
 sky130_fd_sc_hd__nand2_1 _13053_ (.A(_06664_),
    .B(\core.reg_next_pc[8] ),
    .Y(_06774_));
 sky130_fd_sc_hd__a21bo_1 _13054_ (.A1(_06773_),
    .A2(_06662_),
    .B1_N(_06774_),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _13055_ (.A(_06597_),
    .B(\core.reg_out[9] ),
    .Y(_06775_));
 sky130_fd_sc_hd__clkbuf_2 _13056_ (.A(_06620_),
    .X(_06776_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(_06776_),
    .B(\core.alu_out_q[9] ),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_1 _13058_ (.A(_06775_),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_1 _13059_ (.A(_06778_),
    .B(_06008_),
    .Y(_06779_));
 sky130_fd_sc_hd__nand2_1 _13060_ (.A(_05957_),
    .B(\core.reg_next_pc[9] ),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_2 _13061_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__inv_2 _13062_ (.A(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__inv_2 _13063_ (.A(\core.decoded_imm_j[9] ),
    .Y(_06783_));
 sky130_fd_sc_hd__nand2_1 _13064_ (.A(_06782_),
    .B(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__nand2_1 _13065_ (.A(_06781_),
    .B(\core.decoded_imm_j[9] ),
    .Y(_06785_));
 sky130_fd_sc_hd__nand2_1 _13066_ (.A(_06784_),
    .B(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__inv_2 _13067_ (.A(_06786_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(_06765_),
    .B(_06744_),
    .Y(_06788_));
 sky130_fd_sc_hd__nor2_1 _13069_ (.A(_06745_),
    .B(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__nand2_1 _13070_ (.A(_06691_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__nor2_1 _13071_ (.A(_06743_),
    .B(_06764_),
    .Y(_06791_));
 sky130_fd_sc_hd__inv_2 _13072_ (.A(_06763_),
    .Y(_06792_));
 sky130_fd_sc_hd__o21ai_1 _13073_ (.A1(_06741_),
    .A2(_06792_),
    .B1(_06761_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21oi_1 _13074_ (.A1(_06747_),
    .A2(_06791_),
    .B1(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__nand2_1 _13075_ (.A(_06790_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__or2_1 _13076_ (.A(_06787_),
    .B(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__nand2_1 _13077_ (.A(_06795_),
    .B(_06787_),
    .Y(_06797_));
 sky130_fd_sc_hd__nand2_1 _13078_ (.A(_06770_),
    .B(_06782_),
    .Y(_06798_));
 sky130_fd_sc_hd__nor2_2 _13079_ (.A(_06782_),
    .B(_06770_),
    .Y(_06799_));
 sky130_fd_sc_hd__nor2_1 _13080_ (.A(_06632_),
    .B(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__a32o_1 _13081_ (.A1(_06796_),
    .A2(_06632_),
    .A3(_06797_),
    .B1(_06798_),
    .B2(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(_06801_),
    .A1(_06781_),
    .S(_06682_),
    .X(_06802_));
 sky130_fd_sc_hd__nand2_2 _13083_ (.A(_06664_),
    .B(\core.reg_next_pc[9] ),
    .Y(_06803_));
 sky130_fd_sc_hd__a21bo_1 _13084_ (.A1(_06802_),
    .A2(_06662_),
    .B1_N(_06803_),
    .X(_00125_));
 sky130_fd_sc_hd__clkbuf_2 _13085_ (.A(_06667_),
    .X(_06804_));
 sky130_fd_sc_hd__inv_2 _13086_ (.A(\core.reg_out[10] ),
    .Y(_06805_));
 sky130_fd_sc_hd__nand2_1 _13087_ (.A(_06804_),
    .B(\core.alu_out_q[10] ),
    .Y(_06806_));
 sky130_fd_sc_hd__o21ai_1 _13088_ (.A1(_06804_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand2_2 _13089_ (.A(_06807_),
    .B(_06595_),
    .Y(_06808_));
 sky130_fd_sc_hd__nand2_1 _13090_ (.A(_05963_),
    .B(\core.reg_next_pc[10] ),
    .Y(_06809_));
 sky130_fd_sc_hd__nand2_1 _13091_ (.A(_06808_),
    .B(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13092_ (.A(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__or2_1 _13093_ (.A(_06811_),
    .B(_06799_),
    .X(_06812_));
 sky130_fd_sc_hd__nand2_1 _13094_ (.A(_06799_),
    .B(_06811_),
    .Y(_06813_));
 sky130_fd_sc_hd__and2_1 _13095_ (.A(_06813_),
    .B(_06657_),
    .X(_06814_));
 sky130_fd_sc_hd__nand2_1 _13096_ (.A(_06810_),
    .B(\core.decoded_imm_j[10] ),
    .Y(_06815_));
 sky130_fd_sc_hd__inv_2 _13097_ (.A(\core.decoded_imm_j[10] ),
    .Y(_06816_));
 sky130_fd_sc_hd__nand3_4 _13098_ (.A(_06808_),
    .B(_06816_),
    .C(_06809_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_1 _13099_ (.A(_06815_),
    .B(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__nand2_1 _13100_ (.A(_06797_),
    .B(_06785_),
    .Y(_06819_));
 sky130_fd_sc_hd__xnor2_1 _13101_ (.A(_06818_),
    .B(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__a22o_1 _13102_ (.A1(_06812_),
    .A2(_06814_),
    .B1(_06820_),
    .B2(_06731_),
    .X(_06821_));
 sky130_fd_sc_hd__mux2_8 _13103_ (.A0(_06821_),
    .A1(_06811_),
    .S(_06683_),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_4 _13104_ (.A(_06637_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_1 _13105_ (.A(_06822_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__buf_2 _13106_ (.A(_06616_),
    .X(_06825_));
 sky130_fd_sc_hd__nand2_1 _13107_ (.A(_06825_),
    .B(\core.reg_next_pc[10] ),
    .Y(_06826_));
 sky130_fd_sc_hd__nand2_1 _13108_ (.A(_06824_),
    .B(_06826_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _13109_ (.A(\core.reg_out[11] ),
    .Y(_06827_));
 sky130_fd_sc_hd__nand2_1 _13110_ (.A(_06804_),
    .B(\core.alu_out_q[11] ),
    .Y(_06828_));
 sky130_fd_sc_hd__o21ai_1 _13111_ (.A1(_06804_),
    .A2(_06827_),
    .B1(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_06829_),
    .B(_06595_),
    .Y(_06830_));
 sky130_fd_sc_hd__nand2_2 _13113_ (.A(_05963_),
    .B(\core.reg_next_pc[11] ),
    .Y(_06831_));
 sky130_fd_sc_hd__nand2_2 _13114_ (.A(_06830_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(_06832_),
    .B(_04577_),
    .Y(_06833_));
 sky130_fd_sc_hd__nand3b_1 _13116_ (.A_N(\core.decoded_imm_j[11] ),
    .B(_06830_),
    .C(_06831_),
    .Y(_06834_));
 sky130_fd_sc_hd__nand2_1 _13117_ (.A(_06833_),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__inv_2 _13118_ (.A(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nor2_1 _13119_ (.A(_06818_),
    .B(_06786_),
    .Y(_06837_));
 sky130_fd_sc_hd__nand2_1 _13120_ (.A(_06795_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__inv_2 _13121_ (.A(_06817_),
    .Y(_06839_));
 sky130_fd_sc_hd__o21ai_2 _13122_ (.A1(_06785_),
    .A2(_06839_),
    .B1(_06815_),
    .Y(_06840_));
 sky130_fd_sc_hd__inv_2 _13123_ (.A(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__nand2_1 _13124_ (.A(_06838_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__or2_1 _13125_ (.A(_06836_),
    .B(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_06842_),
    .B(_06836_),
    .Y(_06844_));
 sky130_fd_sc_hd__a21o_1 _13127_ (.A1(_06799_),
    .A2(_06811_),
    .B1(_06832_),
    .X(_06845_));
 sky130_fd_sc_hd__nand3_1 _13128_ (.A(_06799_),
    .B(_06811_),
    .C(_06832_),
    .Y(_06846_));
 sky130_fd_sc_hd__and3_1 _13129_ (.A(_06845_),
    .B(_06846_),
    .C(_06657_),
    .X(_06847_));
 sky130_fd_sc_hd__a31o_1 _13130_ (.A1(_06843_),
    .A2(_06703_),
    .A3(_06844_),
    .B1(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__mux2_1 _13131_ (.A0(_06848_),
    .A1(_06832_),
    .S(_06682_),
    .X(_06849_));
 sky130_fd_sc_hd__nand2_1 _13132_ (.A(_06664_),
    .B(\core.reg_next_pc[11] ),
    .Y(_06850_));
 sky130_fd_sc_hd__a21bo_1 _13133_ (.A1(_06849_),
    .A2(_06662_),
    .B1_N(_06850_),
    .X(_00127_));
 sky130_fd_sc_hd__clkbuf_4 _13134_ (.A(_06631_),
    .X(_06851_));
 sky130_fd_sc_hd__inv_2 _13135_ (.A(\core.reg_out[12] ),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_1 _13136_ (.A(_06600_),
    .B(\core.alu_out_q[12] ),
    .Y(_06853_));
 sky130_fd_sc_hd__o21ai_1 _13137_ (.A1(_06600_),
    .A2(_06852_),
    .B1(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand2_1 _13138_ (.A(_06854_),
    .B(_06008_),
    .Y(_06855_));
 sky130_fd_sc_hd__nand2_1 _13139_ (.A(_06001_),
    .B(\core.reg_next_pc[12] ),
    .Y(_06856_));
 sky130_fd_sc_hd__nand2_1 _13140_ (.A(_06855_),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__inv_2 _13141_ (.A(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand2_2 _13142_ (.A(_06846_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__nor2_1 _13143_ (.A(_06858_),
    .B(_06846_),
    .Y(_06860_));
 sky130_fd_sc_hd__nor2_1 _13144_ (.A(_06731_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__nand2_1 _13145_ (.A(_06857_),
    .B(\core.decoded_imm_j[12] ),
    .Y(_06862_));
 sky130_fd_sc_hd__nand3b_1 _13146_ (.A_N(\core.decoded_imm_j[12] ),
    .B(_06855_),
    .C(_06856_),
    .Y(_06863_));
 sky130_fd_sc_hd__nand2_1 _13147_ (.A(_06862_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_06844_),
    .B(_06833_),
    .Y(_06865_));
 sky130_fd_sc_hd__xnor2_1 _13149_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__clkbuf_2 _13150_ (.A(_06632_),
    .X(_06867_));
 sky130_fd_sc_hd__a22o_1 _13151_ (.A1(_06859_),
    .A2(_06861_),
    .B1(_06866_),
    .B2(_06867_),
    .X(_06868_));
 sky130_fd_sc_hd__buf_2 _13152_ (.A(_06631_),
    .X(_06869_));
 sky130_fd_sc_hd__nand2_2 _13153_ (.A(_06868_),
    .B(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__o21ai_4 _13154_ (.A1(_06851_),
    .A2(_06858_),
    .B1(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__clkbuf_4 _13155_ (.A(_06637_),
    .X(_06872_));
 sky130_fd_sc_hd__nand2_8 _13156_ (.A(_06871_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_8 _13157_ (.A(_06825_),
    .B(\core.reg_next_pc[12] ),
    .Y(_06874_));
 sky130_fd_sc_hd__nand2_4 _13158_ (.A(_06873_),
    .B(_06874_),
    .Y(_00128_));
 sky130_fd_sc_hd__buf_6 _13159_ (.A(_06620_),
    .X(_06875_));
 sky130_fd_sc_hd__inv_2 _13160_ (.A(\core.reg_out[13] ),
    .Y(_06876_));
 sky130_fd_sc_hd__nand2_1 _13161_ (.A(_06875_),
    .B(\core.alu_out_q[13] ),
    .Y(_06877_));
 sky130_fd_sc_hd__o21ai_1 _13162_ (.A1(_06875_),
    .A2(_06876_),
    .B1(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__nand2_1 _13163_ (.A(_06878_),
    .B(_06594_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_2 _13164_ (.A(_05962_),
    .B(\core.reg_next_pc[13] ),
    .Y(_06880_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(_06879_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nand2_1 _13166_ (.A(_06881_),
    .B(\core.decoded_imm_j[13] ),
    .Y(_06882_));
 sky130_fd_sc_hd__nand3b_1 _13167_ (.A_N(\core.decoded_imm_j[13] ),
    .B(_06879_),
    .C(_06880_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_2 _13168_ (.A(_06882_),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__inv_2 _13169_ (.A(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__nor2_1 _13170_ (.A(_06864_),
    .B(_06835_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand2_1 _13171_ (.A(_06886_),
    .B(_06837_),
    .Y(_06887_));
 sky130_fd_sc_hd__inv_2 _13172_ (.A(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand2_1 _13173_ (.A(_06795_),
    .B(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__nand2_1 _13174_ (.A(_06840_),
    .B(_06886_),
    .Y(_06890_));
 sky130_fd_sc_hd__inv_2 _13175_ (.A(_06863_),
    .Y(_06891_));
 sky130_fd_sc_hd__o21a_1 _13176_ (.A1(_06833_),
    .A2(_06891_),
    .B1(_06862_),
    .X(_06892_));
 sky130_fd_sc_hd__nand2_1 _13177_ (.A(_06890_),
    .B(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__inv_2 _13178_ (.A(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _13179_ (.A(_06889_),
    .B(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__or2_1 _13180_ (.A(_06885_),
    .B(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__clkbuf_4 _13181_ (.A(_06607_),
    .X(_06897_));
 sky130_fd_sc_hd__nand2_1 _13182_ (.A(_06895_),
    .B(_06885_),
    .Y(_06898_));
 sky130_fd_sc_hd__o21a_1 _13183_ (.A1(_06881_),
    .A2(_06860_),
    .B1(_06658_),
    .X(_06899_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(_06860_),
    .B(_06881_),
    .Y(_06900_));
 sky130_fd_sc_hd__a32o_1 _13185_ (.A1(_06896_),
    .A2(_06897_),
    .A3(_06898_),
    .B1(_06899_),
    .B2(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__and2_1 _13186_ (.A(_06881_),
    .B(_06683_),
    .X(_06902_));
 sky130_fd_sc_hd__a21oi_1 _13187_ (.A1(_06901_),
    .A2(_06660_),
    .B1(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_06825_),
    .B(net135),
    .Y(_06904_));
 sky130_fd_sc_hd__o21ai_1 _13189_ (.A1(_04457_),
    .A2(_06903_),
    .B1(_06904_),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _13190_ (.A(\core.reg_out[14] ),
    .Y(_06905_));
 sky130_fd_sc_hd__nand2_1 _13191_ (.A(_06776_),
    .B(\core.alu_out_q[14] ),
    .Y(_06906_));
 sky130_fd_sc_hd__o21ai_1 _13192_ (.A1(_06600_),
    .A2(_06905_),
    .B1(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand2_1 _13193_ (.A(_06907_),
    .B(_06008_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_1 _13194_ (.A(_06001_),
    .B(\core.reg_next_pc[14] ),
    .Y(_06909_));
 sky130_fd_sc_hd__nand2_2 _13195_ (.A(_06908_),
    .B(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__inv_2 _13196_ (.A(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(_06857_),
    .B(_06881_),
    .Y(_06912_));
 sky130_fd_sc_hd__or2_1 _13198_ (.A(_06912_),
    .B(_06846_),
    .X(_06913_));
 sky130_fd_sc_hd__nand2_1 _13199_ (.A(_06913_),
    .B(_06911_),
    .Y(_06914_));
 sky130_fd_sc_hd__o21a_1 _13200_ (.A1(_06911_),
    .A2(_06913_),
    .B1(_06658_),
    .X(_06915_));
 sky130_fd_sc_hd__nand2_2 _13201_ (.A(_06910_),
    .B(\core.decoded_imm_j[14] ),
    .Y(_06916_));
 sky130_fd_sc_hd__inv_2 _13202_ (.A(\core.decoded_imm_j[14] ),
    .Y(_06917_));
 sky130_fd_sc_hd__nand3_1 _13203_ (.A(_06908_),
    .B(_06917_),
    .C(_06909_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_2 _13204_ (.A(_06916_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__inv_2 _13205_ (.A(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__nand2_1 _13206_ (.A(_06898_),
    .B(_06882_),
    .Y(_06921_));
 sky130_fd_sc_hd__xor2_1 _13207_ (.A(_06920_),
    .B(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__a22o_1 _13208_ (.A1(_06914_),
    .A2(_06915_),
    .B1(_06922_),
    .B2(_06867_),
    .X(_06923_));
 sky130_fd_sc_hd__nand2_1 _13209_ (.A(_06923_),
    .B(_06869_),
    .Y(_06924_));
 sky130_fd_sc_hd__o21ai_1 _13210_ (.A1(_06851_),
    .A2(_06911_),
    .B1(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2_2 _13211_ (.A(_06925_),
    .B(_06872_),
    .Y(_06926_));
 sky130_fd_sc_hd__nand2_2 _13212_ (.A(_06825_),
    .B(\core.reg_next_pc[14] ),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_1 _13213_ (.A(_06926_),
    .B(_06927_),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_2 _13214_ (.A(\core.reg_out[15] ),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(_06776_),
    .B(\core.alu_out_q[15] ),
    .Y(_06929_));
 sky130_fd_sc_hd__o21ai_1 _13216_ (.A1(_06776_),
    .A2(_06928_),
    .B1(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__nand2_1 _13217_ (.A(_06930_),
    .B(_06008_),
    .Y(_06931_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_05957_),
    .B(\core.reg_next_pc[15] ),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_2 _13219_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__nand2_4 _13220_ (.A(_06910_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_2 _13221_ (.A(_06934_),
    .B(_06900_),
    .Y(_06935_));
 sky130_fd_sc_hd__o21ba_1 _13222_ (.A1(_06911_),
    .A2(_06913_),
    .B1_N(_06933_),
    .X(_06936_));
 sky130_fd_sc_hd__nand2_1 _13223_ (.A(_06885_),
    .B(_06920_),
    .Y(_06937_));
 sky130_fd_sc_hd__inv_2 _13224_ (.A(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__nand2_1 _13225_ (.A(_06895_),
    .B(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__inv_2 _13226_ (.A(_06918_),
    .Y(_06940_));
 sky130_fd_sc_hd__o21ai_1 _13227_ (.A1(_06882_),
    .A2(_06940_),
    .B1(_06916_),
    .Y(_06941_));
 sky130_fd_sc_hd__inv_2 _13228_ (.A(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__nand2_1 _13229_ (.A(_06933_),
    .B(\core.decoded_imm_j[15] ),
    .Y(_06943_));
 sky130_fd_sc_hd__nand3_1 _13230_ (.A(_06931_),
    .B(_06296_),
    .C(_06932_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _13231_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand2_1 _13232_ (.A(_06939_),
    .B(_06942_),
    .Y(_06946_));
 sky130_fd_sc_hd__inv_2 _13233_ (.A(_06945_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2_2 _13234_ (.A(_06946_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__buf_2 _13235_ (.A(_06607_),
    .X(_06949_));
 sky130_fd_sc_hd__nand2_1 _13236_ (.A(_06948_),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__a31o_1 _13237_ (.A1(_06939_),
    .A2(_06942_),
    .A3(_06945_),
    .B1(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__o31ai_2 _13238_ (.A1(_06867_),
    .A2(_06935_),
    .A3(_06936_),
    .B1(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand2_1 _13239_ (.A(_06952_),
    .B(_06851_),
    .Y(_06953_));
 sky130_fd_sc_hd__buf_1 _13240_ (.A(_06682_),
    .X(_06954_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13241_ (.A(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__nand2_1 _13242_ (.A(_06933_),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__nand2_1 _13243_ (.A(_06953_),
    .B(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand2_1 _13244_ (.A(_06957_),
    .B(_06872_),
    .Y(_06958_));
 sky130_fd_sc_hd__nand2_1 _13245_ (.A(_06825_),
    .B(\core.reg_next_pc[15] ),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_1 _13246_ (.A(_06958_),
    .B(_06959_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _13247_ (.A(\core.reg_out[16] ),
    .Y(_06960_));
 sky130_fd_sc_hd__nand2_1 _13248_ (.A(_06875_),
    .B(\core.alu_out_q[16] ),
    .Y(_06961_));
 sky130_fd_sc_hd__o21ai_1 _13249_ (.A1(_06776_),
    .A2(_06960_),
    .B1(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand2_2 _13250_ (.A(_06962_),
    .B(_06594_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand2_4 _13251_ (.A(_05957_),
    .B(\core.reg_next_pc[16] ),
    .Y(_06964_));
 sky130_fd_sc_hd__nand2_8 _13252_ (.A(_06963_),
    .B(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__and2_1 _13253_ (.A(_06965_),
    .B(_06954_),
    .X(_06966_));
 sky130_fd_sc_hd__nand2_2 _13254_ (.A(_06965_),
    .B(\core.decoded_imm_j[16] ),
    .Y(_06967_));
 sky130_fd_sc_hd__nand3_4 _13255_ (.A(_06963_),
    .B(_06297_),
    .C(_06964_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand2_2 _13256_ (.A(_06967_),
    .B(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__inv_2 _13257_ (.A(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__nand2_1 _13258_ (.A(_06948_),
    .B(_06943_),
    .Y(_06971_));
 sky130_fd_sc_hd__xor2_1 _13259_ (.A(_06970_),
    .B(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__clkbuf_2 _13260_ (.A(_06632_),
    .X(_06973_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13261_ (.A(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__nand2_1 _13262_ (.A(_06972_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__nor2_2 _13263_ (.A(_06934_),
    .B(_06913_),
    .Y(_06976_));
 sky130_fd_sc_hd__or2_2 _13264_ (.A(_06965_),
    .B(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__nand2_1 _13265_ (.A(_06976_),
    .B(_06965_),
    .Y(_06978_));
 sky130_fd_sc_hd__nand3_1 _13266_ (.A(_06977_),
    .B(_06665_),
    .C(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__a21oi_1 _13267_ (.A1(_06975_),
    .A2(_06979_),
    .B1(_06955_),
    .Y(_06980_));
 sky130_fd_sc_hd__o21ai_1 _13268_ (.A1(_06966_),
    .A2(_06980_),
    .B1(_06823_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand2_1 _13269_ (.A(_06825_),
    .B(\core.reg_next_pc[16] ),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_1 _13270_ (.A(_06981_),
    .B(_06982_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _13271_ (.A(_06754_),
    .B(\core.alu_out_q[17] ),
    .Y(_06983_));
 sky130_fd_sc_hd__o21ai_1 _13272_ (.A1(_06754_),
    .A2(_05955_),
    .B1(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__inv_2 _13273_ (.A(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__o21ai_4 _13274_ (.A1(_06001_),
    .A2(_06985_),
    .B1(_05964_),
    .Y(_06986_));
 sky130_fd_sc_hd__inv_2 _13275_ (.A(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__inv_2 _13276_ (.A(\core.decoded_imm_j[17] ),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_2 _13277_ (.A(_06987_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__nand2_2 _13278_ (.A(_06986_),
    .B(\core.decoded_imm_j[17] ),
    .Y(_06990_));
 sky130_fd_sc_hd__nand2_1 _13279_ (.A(_06989_),
    .B(_06990_),
    .Y(_06991_));
 sky130_fd_sc_hd__inv_2 _13280_ (.A(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__nand2_8 _13281_ (.A(_06947_),
    .B(_06970_),
    .Y(_06993_));
 sky130_fd_sc_hd__nor3_1 _13282_ (.A(_06937_),
    .B(_06993_),
    .C(_06887_),
    .Y(_06994_));
 sky130_fd_sc_hd__nand2_1 _13283_ (.A(_06795_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nor2_1 _13284_ (.A(_06937_),
    .B(_06993_),
    .Y(_06996_));
 sky130_fd_sc_hd__o21a_2 _13285_ (.A1(_06943_),
    .A2(_06969_),
    .B1(_06967_),
    .X(_06997_));
 sky130_fd_sc_hd__nor2_1 _13286_ (.A(_06945_),
    .B(_06969_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand2_2 _13287_ (.A(_06941_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand2_8 _13288_ (.A(_06997_),
    .B(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__a21oi_4 _13289_ (.A1(_06893_),
    .A2(_06996_),
    .B1(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__nand2_2 _13290_ (.A(_06995_),
    .B(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__or2_1 _13291_ (.A(_06992_),
    .B(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(_07002_),
    .B(_06992_),
    .Y(_07004_));
 sky130_fd_sc_hd__and2_1 _13293_ (.A(_07004_),
    .B(_06609_),
    .X(_07005_));
 sky130_fd_sc_hd__nor2_1 _13294_ (.A(_06631_),
    .B(_06987_),
    .Y(_07006_));
 sky130_fd_sc_hd__nand2_1 _13295_ (.A(_06978_),
    .B(_06987_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand2_4 _13296_ (.A(_06986_),
    .B(_06965_),
    .Y(_07008_));
 sky130_fd_sc_hd__nor3_2 _13297_ (.A(_06934_),
    .B(_07008_),
    .C(_06900_),
    .Y(_07009_));
 sky130_fd_sc_hd__inv_2 _13298_ (.A(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__and3_1 _13299_ (.A(_07007_),
    .B(_07010_),
    .C(_04502_),
    .X(_07011_));
 sky130_fd_sc_hd__a211o_1 _13300_ (.A1(_07003_),
    .A2(_07005_),
    .B1(_07006_),
    .C1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__nand2_2 _13301_ (.A(_07012_),
    .B(_06872_),
    .Y(_07013_));
 sky130_fd_sc_hd__clkbuf_4 _13302_ (.A(_06616_),
    .X(_07014_));
 sky130_fd_sc_hd__nand2_1 _13303_ (.A(_07014_),
    .B(\core.reg_next_pc[17] ),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_1 _13304_ (.A(_07013_),
    .B(_07015_),
    .Y(_00133_));
 sky130_fd_sc_hd__nand2_1 _13305_ (.A(_06667_),
    .B(\core.alu_out_q[18] ),
    .Y(_07016_));
 sky130_fd_sc_hd__o21ai_1 _13306_ (.A1(_06875_),
    .A2(_05975_),
    .B1(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__nand2_1 _13307_ (.A(_07017_),
    .B(_06594_),
    .Y(_07018_));
 sky130_fd_sc_hd__nand2_1 _13308_ (.A(_07018_),
    .B(_05976_),
    .Y(_07019_));
 sky130_fd_sc_hd__clkbuf_2 _13309_ (.A(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__or2_1 _13310_ (.A(\core.decoded_imm_j[18] ),
    .B(_07020_),
    .X(_07021_));
 sky130_fd_sc_hd__nand2_1 _13311_ (.A(_07020_),
    .B(\core.decoded_imm_j[18] ),
    .Y(_07022_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(_07021_),
    .B(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand2_1 _13313_ (.A(_07004_),
    .B(_06990_),
    .Y(_07024_));
 sky130_fd_sc_hd__xnor2_1 _13314_ (.A(_07023_),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__and3_1 _13315_ (.A(_06769_),
    .B(_06760_),
    .C(_06781_),
    .X(_07026_));
 sky130_fd_sc_hd__nand2_1 _13316_ (.A(_07026_),
    .B(_06707_),
    .Y(_07027_));
 sky130_fd_sc_hd__and2_1 _13317_ (.A(_05958_),
    .B(\core.reg_next_pc[11] ),
    .X(_07028_));
 sky130_fd_sc_hd__and2_1 _13318_ (.A(_06829_),
    .B(_06009_),
    .X(_07029_));
 sky130_fd_sc_hd__inv_2 _13319_ (.A(_06912_),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_1 _13320_ (.A(_06934_),
    .B(_07008_),
    .Y(_07031_));
 sky130_fd_sc_hd__o2111ai_1 _13321_ (.A1(_07028_),
    .A2(_07029_),
    .B1(_06810_),
    .C1(_07030_),
    .D1(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(_07027_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__xor2_1 _13323_ (.A(_07020_),
    .B(_07033_),
    .X(_07034_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(_07025_),
    .A1(_07034_),
    .S(_06665_),
    .X(_07035_));
 sky130_fd_sc_hd__nand2_1 _13325_ (.A(_07035_),
    .B(_06660_),
    .Y(_07036_));
 sky130_fd_sc_hd__nand2_1 _13326_ (.A(_07020_),
    .B(_06954_),
    .Y(_07037_));
 sky130_fd_sc_hd__nand2_4 _13327_ (.A(_07036_),
    .B(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__nand2_4 _13328_ (.A(_06664_),
    .B(\core.reg_next_pc[18] ),
    .Y(_07039_));
 sky130_fd_sc_hd__a21bo_1 _13329_ (.A1(_07038_),
    .A2(_06662_),
    .B1_N(_07039_),
    .X(_00134_));
 sky130_fd_sc_hd__nand2_1 _13330_ (.A(_06599_),
    .B(\core.alu_out_q[19] ),
    .Y(_07040_));
 sky130_fd_sc_hd__o21ai_1 _13331_ (.A1(_06754_),
    .A2(_05981_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__nand2_1 _13332_ (.A(_07041_),
    .B(_06007_),
    .Y(_07042_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(_07042_),
    .B(_05984_),
    .Y(_07043_));
 sky130_fd_sc_hd__buf_1 _13334_ (.A(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__or2_1 _13335_ (.A(\core.decoded_imm_j[19] ),
    .B(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__nand2_1 _13336_ (.A(_07044_),
    .B(\core.decoded_imm_j[19] ),
    .Y(_07046_));
 sky130_fd_sc_hd__nand2_1 _13337_ (.A(_07045_),
    .B(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__inv_2 _13338_ (.A(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__nor2_2 _13339_ (.A(_07023_),
    .B(_06991_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_07002_),
    .B(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__o21ai_1 _13341_ (.A1(_06990_),
    .A2(_07023_),
    .B1(_07022_),
    .Y(_07051_));
 sky130_fd_sc_hd__inv_2 _13342_ (.A(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(_07050_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__or2_1 _13344_ (.A(_07048_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__nand2_2 _13345_ (.A(_07053_),
    .B(_07048_),
    .Y(_07055_));
 sky130_fd_sc_hd__nand3_1 _13346_ (.A(_07054_),
    .B(_06897_),
    .C(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand2_2 _13347_ (.A(_07033_),
    .B(_07020_),
    .Y(_07057_));
 sky130_fd_sc_hd__or2_1 _13348_ (.A(_07044_),
    .B(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_07057_),
    .B(_07044_),
    .Y(_07059_));
 sky130_fd_sc_hd__a21o_2 _13350_ (.A1(_07058_),
    .A2(_07059_),
    .B1(_06703_),
    .X(_07060_));
 sky130_fd_sc_hd__nand2_1 _13351_ (.A(_07056_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(_07061_),
    .A1(_07044_),
    .S(_06682_),
    .X(_07062_));
 sky130_fd_sc_hd__nand2_8 _13353_ (.A(_06616_),
    .B(\core.reg_next_pc[19] ),
    .Y(_07063_));
 sky130_fd_sc_hd__a21bo_1 _13354_ (.A1(_07062_),
    .A2(_06662_),
    .B1_N(_07063_),
    .X(_00135_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(_07019_),
    .B(_07043_),
    .Y(_07064_));
 sky130_fd_sc_hd__inv_2 _13356_ (.A(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand2_2 _13357_ (.A(_06804_),
    .B(\core.alu_out_q[20] ),
    .Y(_07066_));
 sky130_fd_sc_hd__o21ai_1 _13358_ (.A1(_06804_),
    .A2(_05988_),
    .B1(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__nand2_1 _13359_ (.A(_07067_),
    .B(_06595_),
    .Y(_07068_));
 sky130_fd_sc_hd__nand2_1 _13360_ (.A(_07068_),
    .B(_05991_),
    .Y(_07069_));
 sky130_fd_sc_hd__clkbuf_2 _13361_ (.A(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__a21oi_1 _13362_ (.A1(net104),
    .A2(_07065_),
    .B1(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__nand3_4 _13363_ (.A(net104),
    .B(_07065_),
    .C(_07070_),
    .Y(_07072_));
 sky130_fd_sc_hd__nand2_1 _13364_ (.A(_07072_),
    .B(_06665_),
    .Y(_07073_));
 sky130_fd_sc_hd__or2_1 _13365_ (.A(\core.decoded_imm_j[20] ),
    .B(_07069_),
    .X(_07074_));
 sky130_fd_sc_hd__clkbuf_4 _13366_ (.A(\core.decoded_imm_j[20] ),
    .X(_07075_));
 sky130_fd_sc_hd__nand2_1 _13367_ (.A(_07070_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__nand2_2 _13368_ (.A(_07074_),
    .B(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__nand2_1 _13369_ (.A(_07055_),
    .B(_07046_),
    .Y(_07078_));
 sky130_fd_sc_hd__xnor2_1 _13370_ (.A(_07077_),
    .B(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__clkbuf_4 _13371_ (.A(_06731_),
    .X(_07080_));
 sky130_fd_sc_hd__nand2_1 _13372_ (.A(_07079_),
    .B(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__o21ai_1 _13373_ (.A1(_07071_),
    .A2(_07073_),
    .B1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__nand2_1 _13374_ (.A(_07082_),
    .B(_06851_),
    .Y(_07083_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13375_ (.A(_06954_),
    .X(_07084_));
 sky130_fd_sc_hd__nand2_1 _13376_ (.A(_07070_),
    .B(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__nand2_1 _13377_ (.A(_07083_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(_07086_),
    .B(_06872_),
    .Y(_07087_));
 sky130_fd_sc_hd__nand2_1 _13379_ (.A(_07014_),
    .B(net133),
    .Y(_07088_));
 sky130_fd_sc_hd__nand2_1 _13380_ (.A(_07087_),
    .B(_07088_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_2 _13381_ (.A(_06667_),
    .B(\core.alu_out_q[21] ),
    .Y(_07089_));
 sky130_fd_sc_hd__o21ai_1 _13382_ (.A1(_06667_),
    .A2(_05995_),
    .B1(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__nand2_1 _13383_ (.A(_07090_),
    .B(_06594_),
    .Y(_07091_));
 sky130_fd_sc_hd__nand2_1 _13384_ (.A(_07091_),
    .B(_05996_),
    .Y(_07092_));
 sky130_fd_sc_hd__inv_2 _13385_ (.A(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__nor2_2 _13386_ (.A(_07077_),
    .B(_07047_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_2 _13387_ (.A(_07049_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__inv_2 _13388_ (.A(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__nand2_1 _13389_ (.A(_07002_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__nand2_1 _13390_ (.A(_07051_),
    .B(_07094_),
    .Y(_07098_));
 sky130_fd_sc_hd__o21a_1 _13391_ (.A1(_07046_),
    .A2(_07077_),
    .B1(_07076_),
    .X(_07099_));
 sky130_fd_sc_hd__nand2_4 _13392_ (.A(_07098_),
    .B(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__inv_2 _13393_ (.A(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__inv_2 _13394_ (.A(\core.decoded_imm_j[20] ),
    .Y(_07102_));
 sky130_fd_sc_hd__nand2_2 _13395_ (.A(_07093_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__nand2_2 _13396_ (.A(_07092_),
    .B(\core.decoded_imm_j[20] ),
    .Y(_07104_));
 sky130_fd_sc_hd__nand2_1 _13397_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__nand2_2 _13398_ (.A(_07097_),
    .B(_07101_),
    .Y(_07106_));
 sky130_fd_sc_hd__inv_2 _13399_ (.A(_07105_),
    .Y(_07107_));
 sky130_fd_sc_hd__nand2_1 _13400_ (.A(_07106_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__nand2_4 _13401_ (.A(_07108_),
    .B(_06609_),
    .Y(_07109_));
 sky130_fd_sc_hd__a31o_1 _13402_ (.A1(_07097_),
    .A2(_07101_),
    .A3(_07105_),
    .B1(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__and3_2 _13403_ (.A(_07065_),
    .B(_07070_),
    .C(_07092_),
    .X(_07111_));
 sky130_fd_sc_hd__inv_2 _13404_ (.A(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o21ai_4 _13405_ (.A1(_07112_),
    .A2(_07010_),
    .B1(_04502_),
    .Y(_07113_));
 sky130_fd_sc_hd__a21o_1 _13406_ (.A1(_07072_),
    .A2(_07093_),
    .B1(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__o211ai_2 _13407_ (.A1(_06660_),
    .A2(_07093_),
    .B1(_07110_),
    .C1(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__nand2_1 _13408_ (.A(_07115_),
    .B(_06872_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(_07014_),
    .B(\core.reg_next_pc[21] ),
    .Y(_07117_));
 sky130_fd_sc_hd__nand2_1 _13410_ (.A(_07116_),
    .B(_07117_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _13411_ (.A(_06600_),
    .B(\core.alu_out_q[22] ),
    .Y(_07118_));
 sky130_fd_sc_hd__o21ai_2 _13412_ (.A1(_06600_),
    .A2(_06000_),
    .B1(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__nand2_1 _13413_ (.A(_07119_),
    .B(_06008_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand2_2 _13414_ (.A(_07120_),
    .B(_06002_),
    .Y(_07121_));
 sky130_fd_sc_hd__clkbuf_2 _13415_ (.A(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__and2_1 _13416_ (.A(_07122_),
    .B(_06954_),
    .X(_07123_));
 sky130_fd_sc_hd__or2_1 _13417_ (.A(\core.decoded_imm_j[20] ),
    .B(_07121_),
    .X(_07124_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(_07121_),
    .B(\core.decoded_imm_j[20] ),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_2 _13419_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__inv_2 _13420_ (.A(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_1 _13421_ (.A(_07108_),
    .B(_07104_),
    .Y(_07128_));
 sky130_fd_sc_hd__xor2_1 _13422_ (.A(_07127_),
    .B(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__nand2_1 _13423_ (.A(_07129_),
    .B(_06974_),
    .Y(_07130_));
 sky130_fd_sc_hd__nand2_2 _13424_ (.A(_07033_),
    .B(_07111_),
    .Y(_07131_));
 sky130_fd_sc_hd__or2_1 _13425_ (.A(_07122_),
    .B(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand2_1 _13426_ (.A(_07131_),
    .B(_07122_),
    .Y(_07133_));
 sky130_fd_sc_hd__a21o_1 _13427_ (.A1(_07132_),
    .A2(_07133_),
    .B1(_06867_),
    .X(_07134_));
 sky130_fd_sc_hd__a21oi_1 _13428_ (.A1(_07130_),
    .A2(_07134_),
    .B1(_06955_),
    .Y(_07135_));
 sky130_fd_sc_hd__o21ai_1 _13429_ (.A1(_07123_),
    .A2(_07135_),
    .B1(_06823_),
    .Y(_07136_));
 sky130_fd_sc_hd__nand2_1 _13430_ (.A(_07014_),
    .B(net113),
    .Y(_07137_));
 sky130_fd_sc_hd__nand2_1 _13431_ (.A(_07136_),
    .B(_07137_),
    .Y(_00138_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(\core.reg_out[23] ),
    .A1(\core.alu_out_q[23] ),
    .S(_06667_),
    .X(_07138_));
 sky130_fd_sc_hd__nand2_2 _13433_ (.A(_07138_),
    .B(_06009_),
    .Y(_07139_));
 sky130_fd_sc_hd__nand2_4 _13434_ (.A(_07139_),
    .B(_06012_),
    .Y(_07140_));
 sky130_fd_sc_hd__and2_1 _13435_ (.A(_07140_),
    .B(_06954_),
    .X(_07141_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(_07140_),
    .B(_07075_),
    .Y(_07142_));
 sky130_fd_sc_hd__nand3_2 _13437_ (.A(_07139_),
    .B(_07102_),
    .C(_06012_),
    .Y(_07143_));
 sky130_fd_sc_hd__nand2_1 _13438_ (.A(_07142_),
    .B(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__inv_2 _13439_ (.A(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__nor2_2 _13440_ (.A(_07105_),
    .B(_07126_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand2_1 _13441_ (.A(_07106_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__nand2_1 _13442_ (.A(_07104_),
    .B(_07125_),
    .Y(_07148_));
 sky130_fd_sc_hd__inv_2 _13443_ (.A(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_2 _13444_ (.A(_07147_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_07145_),
    .B(_07150_),
    .X(_07151_));
 sky130_fd_sc_hd__nand2_2 _13446_ (.A(_07150_),
    .B(_07145_),
    .Y(_07152_));
 sky130_fd_sc_hd__nand3_1 _13447_ (.A(_07151_),
    .B(_06974_),
    .C(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__nand2b_1 _13448_ (.A_N(_07131_),
    .B(_07122_),
    .Y(_07154_));
 sky130_fd_sc_hd__or2_1 _13449_ (.A(_07140_),
    .B(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__nand2_1 _13450_ (.A(_07154_),
    .B(_07140_),
    .Y(_07156_));
 sky130_fd_sc_hd__a21o_1 _13451_ (.A1(_07155_),
    .A2(_07156_),
    .B1(_06867_),
    .X(_07157_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(_07153_),
    .A2(_07157_),
    .B1(_06955_),
    .Y(_07158_));
 sky130_fd_sc_hd__o21ai_1 _13453_ (.A1(_07141_),
    .A2(_07158_),
    .B1(_06823_),
    .Y(_07159_));
 sky130_fd_sc_hd__nand2_1 _13454_ (.A(_07014_),
    .B(net116),
    .Y(_07160_));
 sky130_fd_sc_hd__nand2_1 _13455_ (.A(_07159_),
    .B(_07160_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(_07152_),
    .B(_07142_),
    .Y(_07161_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(\core.reg_out[24] ),
    .A1(\core.alu_out_q[24] ),
    .S(_06754_),
    .X(_07162_));
 sky130_fd_sc_hd__nand2_2 _13458_ (.A(_07162_),
    .B(_06595_),
    .Y(_07163_));
 sky130_fd_sc_hd__nand2_2 _13459_ (.A(_07163_),
    .B(_06016_),
    .Y(_07164_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(_07164_),
    .B(_07075_),
    .Y(_07165_));
 sky130_fd_sc_hd__nand3_1 _13461_ (.A(_07163_),
    .B(_07102_),
    .C(_06016_),
    .Y(_07166_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(_07165_),
    .B(_07166_),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_1 _13463_ (.A(_07161_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__inv_2 _13464_ (.A(_07167_),
    .Y(_07169_));
 sky130_fd_sc_hd__nand3_1 _13465_ (.A(_07152_),
    .B(_07142_),
    .C(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(_07168_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2_1 _13467_ (.A(_07171_),
    .B(_07080_),
    .Y(_07172_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_07140_),
    .B(_07122_),
    .Y(_07173_));
 sky130_fd_sc_hd__or2_1 _13469_ (.A(_07173_),
    .B(_07131_),
    .X(_07174_));
 sky130_fd_sc_hd__or2_1 _13470_ (.A(_07164_),
    .B(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__nand2_1 _13471_ (.A(_07174_),
    .B(_07164_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21o_1 _13472_ (.A1(_07175_),
    .A2(_07176_),
    .B1(_06973_),
    .X(_07177_));
 sky130_fd_sc_hd__nand2_1 _13473_ (.A(_07172_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _13474_ (.A(_07178_),
    .B(_06851_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand2_1 _13475_ (.A(_07164_),
    .B(_07084_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _13476_ (.A(_07179_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__buf_2 _13477_ (.A(_06637_),
    .X(_07182_));
 sky130_fd_sc_hd__nand2_1 _13478_ (.A(_07181_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand2_2 _13479_ (.A(_07014_),
    .B(net188),
    .Y(_07184_));
 sky130_fd_sc_hd__nand2_1 _13480_ (.A(_07183_),
    .B(_07184_),
    .Y(_00140_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(\core.reg_out[25] ),
    .A1(\core.alu_out_q[25] ),
    .S(_06875_),
    .X(_07185_));
 sky130_fd_sc_hd__a21oi_4 _13482_ (.A1(_07185_),
    .A2(_06009_),
    .B1(_06023_),
    .Y(_07186_));
 sky130_fd_sc_hd__inv_2 _13483_ (.A(_07164_),
    .Y(_07187_));
 sky130_fd_sc_hd__nor2_1 _13484_ (.A(_07187_),
    .B(_07174_),
    .Y(_07188_));
 sky130_fd_sc_hd__xor2_2 _13485_ (.A(_07186_),
    .B(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__inv_2 _13486_ (.A(_07146_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2_2 _13487_ (.A(_07145_),
    .B(_07169_),
    .Y(_07191_));
 sky130_fd_sc_hd__nor3_1 _13488_ (.A(_07190_),
    .B(_07095_),
    .C(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__nand2_1 _13489_ (.A(_07002_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__nor2_1 _13490_ (.A(_07190_),
    .B(_07191_),
    .Y(_07194_));
 sky130_fd_sc_hd__nand3_2 _13491_ (.A(_07145_),
    .B(_07169_),
    .C(_07148_),
    .Y(_07195_));
 sky130_fd_sc_hd__and2_1 _13492_ (.A(_07142_),
    .B(_07165_),
    .X(_07196_));
 sky130_fd_sc_hd__nand2_1 _13493_ (.A(_07195_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__a21oi_2 _13494_ (.A1(_07100_),
    .A2(_07194_),
    .B1(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__clkinvlp_2 _13495_ (.A(_07186_),
    .Y(_07199_));
 sky130_fd_sc_hd__clkbuf_2 _13496_ (.A(_07075_),
    .X(_07200_));
 sky130_fd_sc_hd__nand2_2 _13497_ (.A(_07199_),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__clkbuf_4 _13498_ (.A(_07102_),
    .X(_07202_));
 sky130_fd_sc_hd__nand2_2 _13499_ (.A(_07186_),
    .B(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__nand2_2 _13500_ (.A(_07201_),
    .B(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_2 _13501_ (.A(_07193_),
    .B(_07198_),
    .Y(_07205_));
 sky130_fd_sc_hd__inv_2 _13502_ (.A(_07204_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_1 _13503_ (.A(_07205_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand2_1 _13504_ (.A(_07207_),
    .B(_06731_),
    .Y(_07208_));
 sky130_fd_sc_hd__a31o_1 _13505_ (.A1(_07193_),
    .A2(_07198_),
    .A3(_07204_),
    .B1(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__o21ai_4 _13506_ (.A1(_07080_),
    .A2(_07189_),
    .B1(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__nand2_1 _13507_ (.A(_07210_),
    .B(_06869_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_1 _13508_ (.A1(_06851_),
    .A2(_07186_),
    .B1(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__nand2_1 _13509_ (.A(_07212_),
    .B(_07182_),
    .Y(_07213_));
 sky130_fd_sc_hd__clkbuf_2 _13510_ (.A(_06616_),
    .X(_07214_));
 sky130_fd_sc_hd__nand2_1 _13511_ (.A(_07214_),
    .B(\core.reg_next_pc[25] ),
    .Y(_07215_));
 sky130_fd_sc_hd__nand2_1 _13512_ (.A(_07213_),
    .B(_07215_),
    .Y(_00141_));
 sky130_fd_sc_hd__mux2_2 _13513_ (.A0(\core.reg_out[26] ),
    .A1(\core.alu_out_q[26] ),
    .S(_06776_),
    .X(_07216_));
 sky130_fd_sc_hd__a21oi_4 _13514_ (.A1(_07216_),
    .A2(_06009_),
    .B1(_06028_),
    .Y(_07217_));
 sky130_fd_sc_hd__nor2_1 _13515_ (.A(_06660_),
    .B(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__inv_2 _13516_ (.A(_07217_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_2 _13517_ (.A(_07219_),
    .B(_07200_),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_1 _13518_ (.A(_07217_),
    .B(_07202_),
    .Y(_07221_));
 sky130_fd_sc_hd__nand2_1 _13519_ (.A(_07220_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__nand2_1 _13520_ (.A(_07207_),
    .B(_07201_),
    .Y(_07223_));
 sky130_fd_sc_hd__xnor2_1 _13521_ (.A(_07222_),
    .B(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__nand2_1 _13522_ (.A(_07224_),
    .B(_06974_),
    .Y(_07225_));
 sky130_fd_sc_hd__or3_2 _13523_ (.A(_07186_),
    .B(_07187_),
    .C(_07173_),
    .X(_07226_));
 sky130_fd_sc_hd__nor3b_4 _13524_ (.A(_07112_),
    .B(_07226_),
    .C_N(_07033_),
    .Y(_07227_));
 sky130_fd_sc_hd__or2_1 _13525_ (.A(_07217_),
    .B(_07227_),
    .X(_07228_));
 sky130_fd_sc_hd__nand2_1 _13526_ (.A(_07227_),
    .B(_07217_),
    .Y(_07229_));
 sky130_fd_sc_hd__a21o_1 _13527_ (.A1(_07228_),
    .A2(_07229_),
    .B1(_06867_),
    .X(_07230_));
 sky130_fd_sc_hd__a21oi_1 _13528_ (.A1(_07225_),
    .A2(_07230_),
    .B1(_06955_),
    .Y(_07231_));
 sky130_fd_sc_hd__o21ai_1 _13529_ (.A1(_07218_),
    .A2(_07231_),
    .B1(_06823_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_1 _13530_ (.A(_07214_),
    .B(\core.reg_next_pc[26] ),
    .Y(_07233_));
 sky130_fd_sc_hd__nand2_1 _13531_ (.A(_07232_),
    .B(_07233_),
    .Y(_00142_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(\core.reg_out[27] ),
    .A1(\core.alu_out_q[27] ),
    .S(_06599_),
    .X(_07234_));
 sky130_fd_sc_hd__a21oi_4 _13533_ (.A1(_07234_),
    .A2(_06595_),
    .B1(_06034_),
    .Y(_07235_));
 sky130_fd_sc_hd__nor2_1 _13534_ (.A(_06660_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__inv_2 _13535_ (.A(_07235_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_4 _13536_ (.A(_07237_),
    .B(_07075_),
    .Y(_07238_));
 sky130_fd_sc_hd__nand2_1 _13537_ (.A(_07235_),
    .B(_07102_),
    .Y(_07239_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(_07238_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__inv_2 _13539_ (.A(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__nor2_1 _13540_ (.A(_07204_),
    .B(_07222_),
    .Y(_07242_));
 sky130_fd_sc_hd__nand2_2 _13541_ (.A(_07205_),
    .B(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__and2_1 _13542_ (.A(_07220_),
    .B(_07201_),
    .X(_07244_));
 sky130_fd_sc_hd__nand2_1 _13543_ (.A(_07243_),
    .B(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__or2_1 _13544_ (.A(_07241_),
    .B(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(_07245_),
    .B(_07241_),
    .Y(_07247_));
 sky130_fd_sc_hd__nand3_1 _13546_ (.A(_07246_),
    .B(_06974_),
    .C(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__nand2_1 _13547_ (.A(_07227_),
    .B(_07219_),
    .Y(_07249_));
 sky130_fd_sc_hd__xor2_1 _13548_ (.A(_07235_),
    .B(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__nand2_1 _13549_ (.A(_07250_),
    .B(_06665_),
    .Y(_07251_));
 sky130_fd_sc_hd__a21oi_1 _13550_ (.A1(_07248_),
    .A2(_07251_),
    .B1(_06955_),
    .Y(_07252_));
 sky130_fd_sc_hd__o21ai_1 _13551_ (.A1(_07236_),
    .A2(_07252_),
    .B1(_06823_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand2_1 _13552_ (.A(_07214_),
    .B(\core.reg_next_pc[27] ),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(_07253_),
    .B(_07254_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _13554_ (.A(_07247_),
    .B(_07238_),
    .Y(_07255_));
 sky130_fd_sc_hd__mux2_2 _13555_ (.A0(\core.reg_out[28] ),
    .A1(\core.alu_out_q[28] ),
    .S(_06875_),
    .X(_07256_));
 sky130_fd_sc_hd__a21oi_2 _13556_ (.A1(_07256_),
    .A2(_06009_),
    .B1(_06040_),
    .Y(_07257_));
 sky130_fd_sc_hd__inv_2 _13557_ (.A(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_07258_),
    .B(_07075_),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_2 _13559_ (.A(_07257_),
    .B(_07102_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_2 _13560_ (.A(_07259_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__nand2_1 _13561_ (.A(_07255_),
    .B(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__inv_2 _13562_ (.A(_07261_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand3_1 _13563_ (.A(_07247_),
    .B(_07238_),
    .C(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__nand2_1 _13564_ (.A(_07262_),
    .B(_07264_),
    .Y(_07265_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(_07265_),
    .B(_07080_),
    .Y(_07266_));
 sky130_fd_sc_hd__buf_4 _13566_ (.A(_07258_),
    .X(_07267_));
 sky130_fd_sc_hd__nand2_2 _13567_ (.A(_07219_),
    .B(_07237_),
    .Y(_07268_));
 sky130_fd_sc_hd__inv_2 _13568_ (.A(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__nand2_1 _13569_ (.A(_07227_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__or2_1 _13570_ (.A(_07267_),
    .B(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__nand2_1 _13571_ (.A(_07270_),
    .B(_07267_),
    .Y(_07272_));
 sky130_fd_sc_hd__a21o_1 _13572_ (.A1(_07271_),
    .A2(_07272_),
    .B1(_06973_),
    .X(_07273_));
 sky130_fd_sc_hd__nand2_1 _13573_ (.A(_07266_),
    .B(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__nand2_4 _13574_ (.A(_07274_),
    .B(_06869_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand2_2 _13575_ (.A(_07267_),
    .B(_07084_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(_07275_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__nand2_1 _13577_ (.A(_07277_),
    .B(_07182_),
    .Y(_07278_));
 sky130_fd_sc_hd__nand2_1 _13578_ (.A(_07214_),
    .B(\core.reg_next_pc[28] ),
    .Y(_07279_));
 sky130_fd_sc_hd__nand2_1 _13579_ (.A(_07278_),
    .B(_07279_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand3b_4 _13580_ (.A_N(_07226_),
    .B(net104),
    .C(_07111_),
    .Y(_07280_));
 sky130_fd_sc_hd__nor2_1 _13581_ (.A(_07268_),
    .B(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__mux2_2 _13582_ (.A0(\core.reg_out[29] ),
    .A1(\core.alu_out_q[29] ),
    .S(_06601_),
    .X(_07282_));
 sky130_fd_sc_hd__a21oi_1 _13583_ (.A1(_07282_),
    .A2(_06010_),
    .B1(_06046_),
    .Y(_07283_));
 sky130_fd_sc_hd__inv_2 _13584_ (.A(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__nand3_4 _13585_ (.A(_07281_),
    .B(_07267_),
    .C(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__inv_2 _13586_ (.A(_07008_),
    .Y(_07286_));
 sky130_fd_sc_hd__nand3_1 _13587_ (.A(_06976_),
    .B(_07286_),
    .C(_07111_),
    .Y(_07287_));
 sky130_fd_sc_hd__nor2_1 _13588_ (.A(_07226_),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand3_4 _13589_ (.A(_07288_),
    .B(_07269_),
    .C(_07267_),
    .Y(_07289_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(_07289_),
    .B(_07283_),
    .Y(_07290_));
 sky130_fd_sc_hd__nand3_1 _13591_ (.A(_07285_),
    .B(_04502_),
    .C(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__and3_1 _13592_ (.A(_07242_),
    .B(_07241_),
    .C(_07263_),
    .X(_07292_));
 sky130_fd_sc_hd__nand2_2 _13593_ (.A(_07205_),
    .B(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__a41o_1 _13594_ (.A1(_07186_),
    .A2(_07217_),
    .A3(_07235_),
    .A4(_07257_),
    .B1(_07202_),
    .X(_07294_));
 sky130_fd_sc_hd__nand2_4 _13595_ (.A(_07284_),
    .B(_07200_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(_07283_),
    .B(_07202_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_2 _13597_ (.A(_07295_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__nand2_2 _13598_ (.A(_07293_),
    .B(_07294_),
    .Y(_07298_));
 sky130_fd_sc_hd__inv_2 _13599_ (.A(_07297_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_2 _13600_ (.A(_07298_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__nand2_4 _13601_ (.A(_07300_),
    .B(_06609_),
    .Y(_07301_));
 sky130_fd_sc_hd__a31o_1 _13602_ (.A1(_07293_),
    .A2(_07294_),
    .A3(_07297_),
    .B1(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__nand2_1 _13603_ (.A(_07284_),
    .B(_07084_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand3_1 _13604_ (.A(_07291_),
    .B(_07302_),
    .C(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__nand2_1 _13605_ (.A(_07304_),
    .B(_07182_),
    .Y(_07305_));
 sky130_fd_sc_hd__nand2_2 _13606_ (.A(_07214_),
    .B(\core.reg_next_pc[29] ),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(_07305_),
    .B(_07306_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand2_2 _13608_ (.A(_07300_),
    .B(_07295_),
    .Y(_07307_));
 sky130_fd_sc_hd__mux2_2 _13609_ (.A0(\core.reg_out[30] ),
    .A1(\core.alu_out_q[30] ),
    .S(_06601_),
    .X(_07308_));
 sky130_fd_sc_hd__a21o_1 _13610_ (.A1(_07308_),
    .A2(_06010_),
    .B1(_06051_),
    .X(_07309_));
 sky130_fd_sc_hd__or2_1 _13611_ (.A(_07200_),
    .B(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__buf_2 _13612_ (.A(_07309_),
    .X(_07311_));
 sky130_fd_sc_hd__nand2_1 _13613_ (.A(_07311_),
    .B(_07200_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_2 _13614_ (.A(_07310_),
    .B(_07312_),
    .Y(_07313_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(_07307_),
    .B(_07313_),
    .Y(_07314_));
 sky130_fd_sc_hd__inv_2 _13616_ (.A(_07313_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand3_2 _13617_ (.A(_07300_),
    .B(_07295_),
    .C(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand2_1 _13618_ (.A(_07314_),
    .B(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__nand2_1 _13619_ (.A(_07317_),
    .B(_07080_),
    .Y(_07318_));
 sky130_fd_sc_hd__and3_1 _13620_ (.A(_07269_),
    .B(_07258_),
    .C(_07284_),
    .X(_07319_));
 sky130_fd_sc_hd__nand2_1 _13621_ (.A(_07227_),
    .B(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__or2_1 _13622_ (.A(_07311_),
    .B(_07320_),
    .X(_07321_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(_07320_),
    .B(_07311_),
    .Y(_07322_));
 sky130_fd_sc_hd__a21o_1 _13624_ (.A1(_07321_),
    .A2(_07322_),
    .B1(_06973_),
    .X(_07323_));
 sky130_fd_sc_hd__nand2_1 _13625_ (.A(_07318_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2_2 _13626_ (.A(_07324_),
    .B(_06869_),
    .Y(_07325_));
 sky130_fd_sc_hd__nand2_1 _13627_ (.A(_07311_),
    .B(_07084_),
    .Y(_07326_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(_07325_),
    .B(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_1 _13629_ (.A(_07327_),
    .B(_07182_),
    .Y(_07328_));
 sky130_fd_sc_hd__nand2_2 _13630_ (.A(_07214_),
    .B(\core.reg_next_pc[30] ),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_1 _13631_ (.A(_07328_),
    .B(_07329_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor2_1 _13632_ (.A(_07297_),
    .B(_07313_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand2_2 _13633_ (.A(_07298_),
    .B(_07330_),
    .Y(_07331_));
 sky130_fd_sc_hd__and2_1 _13634_ (.A(_07295_),
    .B(_07312_),
    .X(_07332_));
 sky130_fd_sc_hd__nand2_4 _13635_ (.A(_07331_),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(\core.reg_out[31] ),
    .A1(\core.alu_out_q[31] ),
    .S(_06601_),
    .X(_07334_));
 sky130_fd_sc_hd__a21bo_1 _13637_ (.A1(_07334_),
    .A2(_06010_),
    .B1_N(_06057_),
    .X(_07335_));
 sky130_fd_sc_hd__xor2_1 _13638_ (.A(_07202_),
    .B(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__nand2_2 _13639_ (.A(_07333_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__inv_2 _13640_ (.A(_07336_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand3_4 _13641_ (.A(_07331_),
    .B(_07332_),
    .C(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand2_2 _13642_ (.A(_07337_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_8 _13643_ (.A(_07340_),
    .B(_07080_),
    .Y(_07341_));
 sky130_fd_sc_hd__and3_1 _13644_ (.A(_07227_),
    .B(_07311_),
    .C(_07319_),
    .X(_07342_));
 sky130_fd_sc_hd__xor2_2 _13645_ (.A(_07335_),
    .B(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__nand2_8 _13646_ (.A(_07343_),
    .B(_06665_),
    .Y(_07344_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_07341_),
    .B(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__nand2_1 _13648_ (.A(_07345_),
    .B(_06869_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(_07335_),
    .B(_07084_),
    .Y(_07347_));
 sky130_fd_sc_hd__nand2_2 _13650_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_8 _13651_ (.A(_07348_),
    .B(_07182_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(_06617_),
    .B(\core.reg_next_pc[31] ),
    .Y(_07350_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(_07349_),
    .B(_07350_),
    .Y(_00147_));
 sky130_fd_sc_hd__a22o_1 _13654_ (.A1(\core.reg_pc[1] ),
    .A2(_06617_),
    .B1(_06606_),
    .B2(_06638_),
    .X(_00148_));
 sky130_fd_sc_hd__buf_2 _13655_ (.A(_06616_),
    .X(_07351_));
 sky130_fd_sc_hd__a22o_1 _13656_ (.A1(\core.reg_pc[2] ),
    .A2(_07351_),
    .B1(_06625_),
    .B2(_06638_),
    .X(_00149_));
 sky130_fd_sc_hd__clkbuf_2 _13657_ (.A(_06637_),
    .X(_07352_));
 sky130_fd_sc_hd__a22o_1 _13658_ (.A1(\core.reg_pc[3] ),
    .A2(_07351_),
    .B1(_06644_),
    .B2(_07352_),
    .X(_00150_));
 sky130_fd_sc_hd__a22o_1 _13659_ (.A1(\core.reg_pc[4] ),
    .A2(_07351_),
    .B1(_06672_),
    .B2(_07352_),
    .X(_00151_));
 sky130_fd_sc_hd__a22o_1 _13660_ (.A1(\core.reg_pc[5] ),
    .A2(_07351_),
    .B1(_06698_),
    .B2(_07352_),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_1 _13661_ (.A1(_05122_),
    .A2(_07351_),
    .B1(_06718_),
    .B2(_07352_),
    .X(_00153_));
 sky130_fd_sc_hd__a22o_1 _13662_ (.A1(\core.reg_pc[7] ),
    .A2(_07351_),
    .B1(_06737_),
    .B2(_07352_),
    .X(_00154_));
 sky130_fd_sc_hd__clkbuf_4 _13663_ (.A(_06615_),
    .X(_07353_));
 sky130_fd_sc_hd__a22o_1 _13664_ (.A1(\core.reg_pc[8] ),
    .A2(_07353_),
    .B1(_06760_),
    .B2(_07352_),
    .X(_00155_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13665_ (.A(_06637_),
    .X(_07354_));
 sky130_fd_sc_hd__a22o_1 _13666_ (.A1(\core.reg_pc[9] ),
    .A2(_07353_),
    .B1(_06781_),
    .B2(_07354_),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_1 _13667_ (.A1(\core.reg_pc[10] ),
    .A2(_07353_),
    .B1(_06811_),
    .B2(_07354_),
    .X(_00157_));
 sky130_fd_sc_hd__a22o_1 _13668_ (.A1(\core.reg_pc[11] ),
    .A2(_07353_),
    .B1(_06832_),
    .B2(_07354_),
    .X(_00158_));
 sky130_fd_sc_hd__a22o_1 _13669_ (.A1(\core.reg_pc[12] ),
    .A2(_07353_),
    .B1(_06857_),
    .B2(_07354_),
    .X(_00159_));
 sky130_fd_sc_hd__a22o_1 _13670_ (.A1(\core.reg_pc[13] ),
    .A2(_07353_),
    .B1(_06881_),
    .B2(_07354_),
    .X(_00160_));
 sky130_fd_sc_hd__clkbuf_4 _13671_ (.A(\core.reg_pc[14] ),
    .X(_07355_));
 sky130_fd_sc_hd__clkbuf_4 _13672_ (.A(_06615_),
    .X(_07356_));
 sky130_fd_sc_hd__a22o_1 _13673_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_06910_),
    .B2(_07354_),
    .X(_00161_));
 sky130_fd_sc_hd__clkbuf_4 _13674_ (.A(_06636_),
    .X(_07357_));
 sky130_fd_sc_hd__a22o_1 _13675_ (.A1(_05275_),
    .A2(_07356_),
    .B1(_06933_),
    .B2(_07357_),
    .X(_00162_));
 sky130_fd_sc_hd__a22o_1 _13676_ (.A1(\core.reg_pc[16] ),
    .A2(_07356_),
    .B1(_06965_),
    .B2(_07357_),
    .X(_00163_));
 sky130_fd_sc_hd__a22o_1 _13677_ (.A1(\core.reg_pc[17] ),
    .A2(_07356_),
    .B1(_06986_),
    .B2(_07357_),
    .X(_00164_));
 sky130_fd_sc_hd__a22o_1 _13678_ (.A1(_05339_),
    .A2(_07356_),
    .B1(_07020_),
    .B2(_07357_),
    .X(_00165_));
 sky130_fd_sc_hd__a22o_1 _13679_ (.A1(\core.reg_pc[19] ),
    .A2(_07356_),
    .B1(_07044_),
    .B2(_07357_),
    .X(_00166_));
 sky130_fd_sc_hd__buf_2 _13680_ (.A(_06615_),
    .X(_07358_));
 sky130_fd_sc_hd__a22o_1 _13681_ (.A1(\core.reg_pc[20] ),
    .A2(_07358_),
    .B1(_07070_),
    .B2(_07357_),
    .X(_00167_));
 sky130_fd_sc_hd__buf_2 _13682_ (.A(_06636_),
    .X(_07359_));
 sky130_fd_sc_hd__a22o_1 _13683_ (.A1(\core.reg_pc[21] ),
    .A2(_07358_),
    .B1(_07092_),
    .B2(_07359_),
    .X(_00168_));
 sky130_fd_sc_hd__a22o_1 _13684_ (.A1(\core.reg_pc[22] ),
    .A2(_07358_),
    .B1(_07122_),
    .B2(_07359_),
    .X(_00169_));
 sky130_fd_sc_hd__a22o_1 _13685_ (.A1(\core.reg_pc[23] ),
    .A2(_07358_),
    .B1(_07140_),
    .B2(_07359_),
    .X(_00170_));
 sky130_fd_sc_hd__a22o_1 _13686_ (.A1(\core.reg_pc[24] ),
    .A2(_07358_),
    .B1(_07164_),
    .B2(_07359_),
    .X(_00171_));
 sky130_fd_sc_hd__a22o_1 _13687_ (.A1(\core.reg_pc[25] ),
    .A2(_07358_),
    .B1(_07199_),
    .B2(_07359_),
    .X(_00172_));
 sky130_fd_sc_hd__buf_2 _13688_ (.A(_06615_),
    .X(_07360_));
 sky130_fd_sc_hd__a22o_1 _13689_ (.A1(_05464_),
    .A2(_07360_),
    .B1(_07219_),
    .B2(_07359_),
    .X(_00173_));
 sky130_fd_sc_hd__a22o_1 _13690_ (.A1(\core.reg_pc[27] ),
    .A2(_07360_),
    .B1(_07237_),
    .B2(_06685_),
    .X(_00174_));
 sky130_fd_sc_hd__a22o_1 _13691_ (.A1(_05492_),
    .A2(_07360_),
    .B1(_07267_),
    .B2(_06685_),
    .X(_00175_));
 sky130_fd_sc_hd__a22o_1 _13692_ (.A1(\core.reg_pc[29] ),
    .A2(_07360_),
    .B1(_07284_),
    .B2(_06685_),
    .X(_00176_));
 sky130_fd_sc_hd__a22o_1 _13693_ (.A1(\core.reg_pc[30] ),
    .A2(_07360_),
    .B1(_07311_),
    .B2(_06685_),
    .X(_00177_));
 sky130_fd_sc_hd__a22o_1 _13694_ (.A1(\core.reg_pc[31] ),
    .A2(_07360_),
    .B1(_07335_),
    .B2(_06685_),
    .X(_00178_));
 sky130_fd_sc_hd__nand2_1 _13695_ (.A(\core.cpu_state[1] ),
    .B(\core.decoder_trigger ),
    .Y(_07361_));
 sky130_fd_sc_hd__inv_2 _13696_ (.A(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__buf_1 _13697_ (.A(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__or2_1 _13698_ (.A(\core.count_instr[0] ),
    .B(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__nand2_1 _13699_ (.A(_07363_),
    .B(\core.count_instr[0] ),
    .Y(_07365_));
 sky130_fd_sc_hd__and3_1 _13700_ (.A(_07364_),
    .B(_06451_),
    .C(_07365_),
    .X(_07366_));
 sky130_fd_sc_hd__buf_1 _13701_ (.A(_07366_),
    .X(_00179_));
 sky130_fd_sc_hd__inv_2 _13702_ (.A(\core.count_instr[1] ),
    .Y(_07367_));
 sky130_fd_sc_hd__or2_1 _13703_ (.A(_07367_),
    .B(_07365_),
    .X(_07368_));
 sky130_fd_sc_hd__clkbuf_2 _13704_ (.A(_06357_),
    .X(_07369_));
 sky130_fd_sc_hd__nand2_1 _13705_ (.A(_07365_),
    .B(_07367_),
    .Y(_07370_));
 sky130_fd_sc_hd__and3_1 _13706_ (.A(_07368_),
    .B(_07369_),
    .C(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__buf_1 _13707_ (.A(_07371_),
    .X(_00180_));
 sky130_fd_sc_hd__or2_1 _13708_ (.A(\core.count_instr[2] ),
    .B(_07368_),
    .X(_07372_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(_07368_),
    .B(\core.count_instr[2] ),
    .Y(_07373_));
 sky130_fd_sc_hd__a21oi_1 _13710_ (.A1(_07372_),
    .A2(_07373_),
    .B1(_06582_),
    .Y(_00181_));
 sky130_fd_sc_hd__and3_1 _13711_ (.A(\core.count_instr[2] ),
    .B(\core.count_instr[1] ),
    .C(\core.count_instr[0] ),
    .X(_07374_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13712_ (.A(_07363_),
    .X(_07375_));
 sky130_fd_sc_hd__inv_2 _13713_ (.A(\core.count_instr[3] ),
    .Y(_07376_));
 sky130_fd_sc_hd__a21oi_1 _13714_ (.A1(_07374_),
    .A2(_07375_),
    .B1(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__and3_1 _13715_ (.A(_07374_),
    .B(_07376_),
    .C(_07375_),
    .X(_07378_));
 sky130_fd_sc_hd__o21a_1 _13716_ (.A1(_07377_),
    .A2(_07378_),
    .B1(_06506_),
    .X(_00182_));
 sky130_fd_sc_hd__buf_2 _13717_ (.A(_07361_),
    .X(_07379_));
 sky130_fd_sc_hd__nand2_1 _13718_ (.A(_07374_),
    .B(\core.count_instr[3] ),
    .Y(_07380_));
 sky130_fd_sc_hd__nor2_1 _13719_ (.A(_07379_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__or2_1 _13720_ (.A(\core.count_instr[4] ),
    .B(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__nand2_1 _13721_ (.A(_07381_),
    .B(\core.count_instr[4] ),
    .Y(_07383_));
 sky130_fd_sc_hd__and3_1 _13722_ (.A(_07382_),
    .B(_07369_),
    .C(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__buf_1 _13723_ (.A(_07384_),
    .X(_00183_));
 sky130_fd_sc_hd__or2_1 _13724_ (.A(\core.count_instr[5] ),
    .B(_07383_),
    .X(_07385_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(_07383_),
    .B(\core.count_instr[5] ),
    .Y(_07386_));
 sky130_fd_sc_hd__buf_2 _13726_ (.A(_06520_),
    .X(_07387_));
 sky130_fd_sc_hd__a21oi_1 _13727_ (.A1(_07385_),
    .A2(_07386_),
    .B1(_07387_),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _13728_ (.A(\core.count_instr[6] ),
    .Y(_07388_));
 sky130_fd_sc_hd__nand2_1 _13729_ (.A(\core.count_instr[5] ),
    .B(\core.count_instr[4] ),
    .Y(_07389_));
 sky130_fd_sc_hd__or2_2 _13730_ (.A(_07389_),
    .B(_07380_),
    .X(_07390_));
 sky130_fd_sc_hd__inv_2 _13731_ (.A(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(_07391_),
    .B(_07363_),
    .Y(_07392_));
 sky130_fd_sc_hd__nor2_1 _13733_ (.A(_07388_),
    .B(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__inv_2 _13734_ (.A(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__nand2_1 _13735_ (.A(_07392_),
    .B(_07388_),
    .Y(_07395_));
 sky130_fd_sc_hd__and3_1 _13736_ (.A(_07394_),
    .B(_07369_),
    .C(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__clkbuf_1 _13737_ (.A(_07396_),
    .X(_00185_));
 sky130_fd_sc_hd__or2_1 _13738_ (.A(\core.count_instr[7] ),
    .B(_07394_),
    .X(_07397_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(_07394_),
    .B(\core.count_instr[7] ),
    .Y(_07398_));
 sky130_fd_sc_hd__a21oi_1 _13740_ (.A1(_07397_),
    .A2(_07398_),
    .B1(_07387_),
    .Y(_00186_));
 sky130_fd_sc_hd__and3_2 _13741_ (.A(_07391_),
    .B(\core.count_instr[7] ),
    .C(\core.count_instr[6] ),
    .X(_07399_));
 sky130_fd_sc_hd__inv_2 _13742_ (.A(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__nor2_1 _13743_ (.A(_07379_),
    .B(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__or2_1 _13744_ (.A(\core.count_instr[8] ),
    .B(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__nand2_1 _13745_ (.A(_07401_),
    .B(\core.count_instr[8] ),
    .Y(_07403_));
 sky130_fd_sc_hd__and3_1 _13746_ (.A(_07402_),
    .B(_07369_),
    .C(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__buf_1 _13747_ (.A(_07404_),
    .X(_00187_));
 sky130_fd_sc_hd__or2_1 _13748_ (.A(\core.count_instr[9] ),
    .B(_07403_),
    .X(_07405_));
 sky130_fd_sc_hd__nand2_1 _13749_ (.A(_07403_),
    .B(\core.count_instr[9] ),
    .Y(_07406_));
 sky130_fd_sc_hd__a21oi_1 _13750_ (.A1(_07405_),
    .A2(_07406_),
    .B1(_07387_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _13751_ (.A(\core.count_instr[9] ),
    .B(\core.count_instr[8] ),
    .Y(_07407_));
 sky130_fd_sc_hd__inv_2 _13752_ (.A(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__a31o_1 _13753_ (.A1(_07399_),
    .A2(_07363_),
    .A3(_07408_),
    .B1(\core.count_instr[10] ),
    .X(_07409_));
 sky130_fd_sc_hd__nand3_1 _13754_ (.A(_07401_),
    .B(\core.count_instr[10] ),
    .C(_07408_),
    .Y(_07410_));
 sky130_fd_sc_hd__and3_1 _13755_ (.A(_07409_),
    .B(_07369_),
    .C(_07410_),
    .X(_07411_));
 sky130_fd_sc_hd__buf_1 _13756_ (.A(_07411_),
    .X(_00189_));
 sky130_fd_sc_hd__or2_1 _13757_ (.A(\core.count_instr[11] ),
    .B(_07410_),
    .X(_07412_));
 sky130_fd_sc_hd__nand2_1 _13758_ (.A(_07410_),
    .B(\core.count_instr[11] ),
    .Y(_07413_));
 sky130_fd_sc_hd__a21oi_1 _13759_ (.A1(_07412_),
    .A2(_07413_),
    .B1(_07387_),
    .Y(_00190_));
 sky130_fd_sc_hd__buf_2 _13760_ (.A(_07362_),
    .X(_07414_));
 sky130_fd_sc_hd__and3_1 _13761_ (.A(_07408_),
    .B(\core.count_instr[11] ),
    .C(\core.count_instr[10] ),
    .X(_07415_));
 sky130_fd_sc_hd__and3_1 _13762_ (.A(_07399_),
    .B(_07414_),
    .C(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__or2_1 _13763_ (.A(\core.count_instr[12] ),
    .B(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__nand2_1 _13764_ (.A(_07416_),
    .B(\core.count_instr[12] ),
    .Y(_07418_));
 sky130_fd_sc_hd__and3_1 _13765_ (.A(_07417_),
    .B(_07369_),
    .C(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__buf_1 _13766_ (.A(_07419_),
    .X(_00191_));
 sky130_fd_sc_hd__or2_1 _13767_ (.A(\core.count_instr[13] ),
    .B(_07418_),
    .X(_07420_));
 sky130_fd_sc_hd__nand2_1 _13768_ (.A(_07418_),
    .B(\core.count_instr[13] ),
    .Y(_07421_));
 sky130_fd_sc_hd__a21oi_1 _13769_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_07387_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _13770_ (.A(\core.count_instr[13] ),
    .B(\core.count_instr[12] ),
    .Y(_07422_));
 sky130_fd_sc_hd__inv_2 _13771_ (.A(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__and2_1 _13772_ (.A(_07416_),
    .B(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__or2_1 _13773_ (.A(\core.count_instr[14] ),
    .B(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__buf_1 _13774_ (.A(_06357_),
    .X(_07426_));
 sky130_fd_sc_hd__nand2_1 _13775_ (.A(_07424_),
    .B(\core.count_instr[14] ),
    .Y(_07427_));
 sky130_fd_sc_hd__and3_1 _13776_ (.A(_07425_),
    .B(_07426_),
    .C(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__clkbuf_1 _13777_ (.A(_07428_),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _13778_ (.A(\core.count_instr[15] ),
    .B(_07427_),
    .X(_07429_));
 sky130_fd_sc_hd__nand2_1 _13779_ (.A(_07427_),
    .B(\core.count_instr[15] ),
    .Y(_07430_));
 sky130_fd_sc_hd__a21oi_1 _13780_ (.A1(_07429_),
    .A2(_07430_),
    .B1(_07387_),
    .Y(_00194_));
 sky130_fd_sc_hd__and3_1 _13781_ (.A(_07423_),
    .B(\core.count_instr[15] ),
    .C(\core.count_instr[14] ),
    .X(_07431_));
 sky130_fd_sc_hd__and4_1 _13782_ (.A(_07399_),
    .B(_07414_),
    .C(_07415_),
    .D(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__or2_1 _13783_ (.A(\core.count_instr[16] ),
    .B(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(_07432_),
    .B(\core.count_instr[16] ),
    .Y(_07434_));
 sky130_fd_sc_hd__and3_1 _13785_ (.A(_07433_),
    .B(_07426_),
    .C(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__buf_1 _13786_ (.A(_07435_),
    .X(_00195_));
 sky130_fd_sc_hd__or2_1 _13787_ (.A(\core.count_instr[17] ),
    .B(_07434_),
    .X(_07436_));
 sky130_fd_sc_hd__nand2_1 _13788_ (.A(_07434_),
    .B(\core.count_instr[17] ),
    .Y(_07437_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13789_ (.A(_06520_),
    .X(_07438_));
 sky130_fd_sc_hd__a21oi_1 _13790_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07438_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(\core.count_instr[17] ),
    .B(\core.count_instr[16] ),
    .Y(_07439_));
 sky130_fd_sc_hd__inv_2 _13792_ (.A(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__and2_1 _13793_ (.A(_07432_),
    .B(_07440_),
    .X(_07441_));
 sky130_fd_sc_hd__or2_1 _13794_ (.A(\core.count_instr[18] ),
    .B(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__nand2_2 _13795_ (.A(_07441_),
    .B(\core.count_instr[18] ),
    .Y(_07443_));
 sky130_fd_sc_hd__and3_1 _13796_ (.A(_07442_),
    .B(_07426_),
    .C(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__buf_1 _13797_ (.A(_07444_),
    .X(_00197_));
 sky130_fd_sc_hd__or2_1 _13798_ (.A(\core.count_instr[19] ),
    .B(_07443_),
    .X(_07445_));
 sky130_fd_sc_hd__nand2_1 _13799_ (.A(_07443_),
    .B(\core.count_instr[19] ),
    .Y(_07446_));
 sky130_fd_sc_hd__a21oi_1 _13800_ (.A1(_07445_),
    .A2(_07446_),
    .B1(_07438_),
    .Y(_00198_));
 sky130_fd_sc_hd__and3_2 _13801_ (.A(_07399_),
    .B(_07415_),
    .C(_07431_),
    .X(_07447_));
 sky130_fd_sc_hd__and3_2 _13802_ (.A(_07440_),
    .B(\core.count_instr[19] ),
    .C(\core.count_instr[18] ),
    .X(_07448_));
 sky130_fd_sc_hd__nand2_1 _13803_ (.A(_07447_),
    .B(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__inv_2 _13804_ (.A(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__nand2_1 _13805_ (.A(_07450_),
    .B(_07362_),
    .Y(_07451_));
 sky130_fd_sc_hd__inv_2 _13806_ (.A(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__or2_1 _13807_ (.A(\core.count_instr[20] ),
    .B(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(_07452_),
    .B(\core.count_instr[20] ),
    .Y(_07454_));
 sky130_fd_sc_hd__and3_1 _13809_ (.A(_07453_),
    .B(_07426_),
    .C(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__clkbuf_1 _13810_ (.A(_07455_),
    .X(_00199_));
 sky130_fd_sc_hd__or2_1 _13811_ (.A(\core.count_instr[21] ),
    .B(_07454_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_1 _13812_ (.A(_07454_),
    .B(\core.count_instr[21] ),
    .Y(_07457_));
 sky130_fd_sc_hd__a21oi_1 _13813_ (.A1(_07456_),
    .A2(_07457_),
    .B1(_07438_),
    .Y(_00200_));
 sky130_fd_sc_hd__and3_1 _13814_ (.A(_07452_),
    .B(\core.count_instr[21] ),
    .C(\core.count_instr[20] ),
    .X(_07458_));
 sky130_fd_sc_hd__or2_1 _13815_ (.A(\core.count_instr[22] ),
    .B(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__nand2_1 _13816_ (.A(_07458_),
    .B(\core.count_instr[22] ),
    .Y(_07460_));
 sky130_fd_sc_hd__and3_1 _13817_ (.A(_07459_),
    .B(_07426_),
    .C(_07460_),
    .X(_07461_));
 sky130_fd_sc_hd__clkbuf_1 _13818_ (.A(_07461_),
    .X(_00201_));
 sky130_fd_sc_hd__or2_1 _13819_ (.A(\core.count_instr[23] ),
    .B(_07460_),
    .X(_07462_));
 sky130_fd_sc_hd__nand2_1 _13820_ (.A(_07460_),
    .B(\core.count_instr[23] ),
    .Y(_07463_));
 sky130_fd_sc_hd__a21oi_1 _13821_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07438_),
    .Y(_00202_));
 sky130_fd_sc_hd__and4_1 _13822_ (.A(\core.count_instr[23] ),
    .B(\core.count_instr[22] ),
    .C(\core.count_instr[21] ),
    .D(\core.count_instr[20] ),
    .X(_07464_));
 sky130_fd_sc_hd__nand2_2 _13823_ (.A(_07450_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor2_1 _13824_ (.A(_07361_),
    .B(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__or2_1 _13825_ (.A(\core.count_instr[24] ),
    .B(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(_07466_),
    .B(\core.count_instr[24] ),
    .Y(_07468_));
 sky130_fd_sc_hd__and3_1 _13827_ (.A(_07467_),
    .B(_07426_),
    .C(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__buf_1 _13828_ (.A(_07469_),
    .X(_00203_));
 sky130_fd_sc_hd__or2_1 _13829_ (.A(\core.count_instr[25] ),
    .B(_07468_),
    .X(_07470_));
 sky130_fd_sc_hd__nand2_1 _13830_ (.A(_07468_),
    .B(\core.count_instr[25] ),
    .Y(_07471_));
 sky130_fd_sc_hd__a21oi_1 _13831_ (.A1(_07470_),
    .A2(_07471_),
    .B1(_07438_),
    .Y(_00204_));
 sky130_fd_sc_hd__and3_1 _13832_ (.A(_07466_),
    .B(\core.count_instr[25] ),
    .C(\core.count_instr[24] ),
    .X(_07472_));
 sky130_fd_sc_hd__or2_1 _13833_ (.A(\core.count_instr[26] ),
    .B(_07472_),
    .X(_07473_));
 sky130_fd_sc_hd__clkbuf_2 _13834_ (.A(_06357_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_1 _13835_ (.A(_07472_),
    .B(\core.count_instr[26] ),
    .Y(_07475_));
 sky130_fd_sc_hd__and3_1 _13836_ (.A(_07473_),
    .B(_07474_),
    .C(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__clkbuf_1 _13837_ (.A(_07476_),
    .X(_00205_));
 sky130_fd_sc_hd__or2_1 _13838_ (.A(\core.count_instr[27] ),
    .B(_07475_),
    .X(_07477_));
 sky130_fd_sc_hd__nand2_1 _13839_ (.A(_07475_),
    .B(\core.count_instr[27] ),
    .Y(_07478_));
 sky130_fd_sc_hd__a21oi_1 _13840_ (.A1(_07477_),
    .A2(_07478_),
    .B1(_07438_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _13841_ (.A(\core.count_instr[25] ),
    .B(\core.count_instr[24] ),
    .Y(_07479_));
 sky130_fd_sc_hd__nand2_1 _13842_ (.A(\core.count_instr[27] ),
    .B(\core.count_instr[26] ),
    .Y(_07480_));
 sky130_fd_sc_hd__nor2_2 _13843_ (.A(_07479_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__and3_1 _13844_ (.A(_07450_),
    .B(_07464_),
    .C(_07481_),
    .X(_07482_));
 sky130_fd_sc_hd__nand2_1 _13845_ (.A(_07482_),
    .B(_07414_),
    .Y(_07483_));
 sky130_fd_sc_hd__inv_2 _13846_ (.A(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__or2_1 _13847_ (.A(\core.count_instr[28] ),
    .B(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(_07484_),
    .B(\core.count_instr[28] ),
    .Y(_07486_));
 sky130_fd_sc_hd__and3_1 _13849_ (.A(_07485_),
    .B(_07474_),
    .C(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__buf_1 _13850_ (.A(_07487_),
    .X(_00207_));
 sky130_fd_sc_hd__or2_1 _13851_ (.A(\core.count_instr[29] ),
    .B(_07486_),
    .X(_07488_));
 sky130_fd_sc_hd__nand2_1 _13852_ (.A(_07486_),
    .B(\core.count_instr[29] ),
    .Y(_07489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13853_ (.A(_06520_),
    .X(_07490_));
 sky130_fd_sc_hd__a21oi_1 _13854_ (.A1(_07488_),
    .A2(_07489_),
    .B1(_07490_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(\core.count_instr[29] ),
    .B(\core.count_instr[28] ),
    .Y(_07491_));
 sky130_fd_sc_hd__nor2_2 _13856_ (.A(_07491_),
    .B(_07483_),
    .Y(_07492_));
 sky130_fd_sc_hd__inv_2 _13857_ (.A(_07491_),
    .Y(_07493_));
 sky130_fd_sc_hd__a31o_1 _13858_ (.A1(_07484_),
    .A2(\core.count_instr[30] ),
    .A3(_07493_),
    .B1(_04513_),
    .X(_07494_));
 sky130_fd_sc_hd__o21ba_1 _13859_ (.A1(\core.count_instr[30] ),
    .A2(_07492_),
    .B1_N(_07494_),
    .X(_07495_));
 sky130_fd_sc_hd__clkbuf_1 _13860_ (.A(_07495_),
    .X(_00209_));
 sky130_fd_sc_hd__a21bo_1 _13861_ (.A1(_07492_),
    .A2(\core.count_instr[30] ),
    .B1_N(\core.count_instr[31] ),
    .X(_07496_));
 sky130_fd_sc_hd__nand3b_1 _13862_ (.A_N(\core.count_instr[31] ),
    .B(_07492_),
    .C(\core.count_instr[30] ),
    .Y(_07497_));
 sky130_fd_sc_hd__a21oi_1 _13863_ (.A1(_07496_),
    .A2(_07497_),
    .B1(_07490_),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _13864_ (.A(\core.count_instr[32] ),
    .Y(_07498_));
 sky130_fd_sc_hd__and3_1 _13865_ (.A(_07493_),
    .B(\core.count_instr[31] ),
    .C(\core.count_instr[30] ),
    .X(_07499_));
 sky130_fd_sc_hd__and4_1 _13866_ (.A(_07464_),
    .B(_07448_),
    .C(_07499_),
    .D(_07481_),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_2 _13867_ (.A(_07447_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__nor2_1 _13868_ (.A(_07361_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__inv_2 _13869_ (.A(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__nor2_1 _13870_ (.A(_07498_),
    .B(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__inv_2 _13871_ (.A(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_07503_),
    .B(_07498_),
    .Y(_07506_));
 sky130_fd_sc_hd__and3_2 _13873_ (.A(_07505_),
    .B(_07474_),
    .C(_07506_),
    .X(_07507_));
 sky130_fd_sc_hd__buf_1 _13874_ (.A(_07507_),
    .X(_00211_));
 sky130_fd_sc_hd__nand2_1 _13875_ (.A(_07505_),
    .B(\core.count_instr[33] ),
    .Y(_07508_));
 sky130_fd_sc_hd__inv_2 _13876_ (.A(\core.count_instr[33] ),
    .Y(_07509_));
 sky130_fd_sc_hd__nand2_1 _13877_ (.A(_07504_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__a21oi_1 _13878_ (.A1(_07508_),
    .A2(_07510_),
    .B1(_07490_),
    .Y(_00212_));
 sky130_fd_sc_hd__and3_1 _13879_ (.A(_07502_),
    .B(\core.count_instr[33] ),
    .C(\core.count_instr[32] ),
    .X(_07511_));
 sky130_fd_sc_hd__or2_1 _13880_ (.A(\core.count_instr[34] ),
    .B(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__nand2_1 _13881_ (.A(_07511_),
    .B(\core.count_instr[34] ),
    .Y(_07513_));
 sky130_fd_sc_hd__and3_1 _13882_ (.A(_07512_),
    .B(_07474_),
    .C(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__buf_1 _13883_ (.A(_07514_),
    .X(_00213_));
 sky130_fd_sc_hd__or2_1 _13884_ (.A(\core.count_instr[35] ),
    .B(_07513_),
    .X(_07515_));
 sky130_fd_sc_hd__nand2_1 _13885_ (.A(_07513_),
    .B(\core.count_instr[35] ),
    .Y(_07516_));
 sky130_fd_sc_hd__a21oi_1 _13886_ (.A1(_07515_),
    .A2(_07516_),
    .B1(_07490_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _13887_ (.A(\core.count_instr[35] ),
    .B(\core.count_instr[34] ),
    .Y(_07517_));
 sky130_fd_sc_hd__or3_2 _13888_ (.A(_07509_),
    .B(_07498_),
    .C(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__nor2_1 _13889_ (.A(_07518_),
    .B(_07501_),
    .Y(_07519_));
 sky130_fd_sc_hd__nand2_1 _13890_ (.A(_07519_),
    .B(_07414_),
    .Y(_07520_));
 sky130_fd_sc_hd__inv_2 _13891_ (.A(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__or2_1 _13892_ (.A(\core.count_instr[36] ),
    .B(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__nand2_1 _13893_ (.A(_07521_),
    .B(\core.count_instr[36] ),
    .Y(_07523_));
 sky130_fd_sc_hd__and3_1 _13894_ (.A(_07522_),
    .B(_07474_),
    .C(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__clkbuf_1 _13895_ (.A(_07524_),
    .X(_00215_));
 sky130_fd_sc_hd__or2_1 _13896_ (.A(\core.count_instr[37] ),
    .B(_07523_),
    .X(_07525_));
 sky130_fd_sc_hd__nand2_1 _13897_ (.A(_07523_),
    .B(\core.count_instr[37] ),
    .Y(_07526_));
 sky130_fd_sc_hd__a21oi_1 _13898_ (.A1(_07525_),
    .A2(_07526_),
    .B1(_07490_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _13899_ (.A(\core.count_instr[38] ),
    .Y(_07527_));
 sky130_fd_sc_hd__nand2_1 _13900_ (.A(\core.count_instr[37] ),
    .B(\core.count_instr[36] ),
    .Y(_07528_));
 sky130_fd_sc_hd__nor2_1 _13901_ (.A(_07528_),
    .B(_07520_),
    .Y(_07529_));
 sky130_fd_sc_hd__inv_2 _13902_ (.A(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__nor2_1 _13903_ (.A(_07527_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__inv_2 _13904_ (.A(_07531_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand2_1 _13905_ (.A(_07530_),
    .B(_07527_),
    .Y(_07533_));
 sky130_fd_sc_hd__and3_1 _13906_ (.A(_07532_),
    .B(_07474_),
    .C(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__buf_1 _13907_ (.A(_07534_),
    .X(_00217_));
 sky130_fd_sc_hd__nand2_1 _13908_ (.A(_07532_),
    .B(\core.count_instr[39] ),
    .Y(_07535_));
 sky130_fd_sc_hd__inv_2 _13909_ (.A(\core.count_instr[39] ),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(_07531_),
    .B(_07536_),
    .Y(_07537_));
 sky130_fd_sc_hd__a21oi_1 _13911_ (.A1(_07535_),
    .A2(_07537_),
    .B1(_07490_),
    .Y(_00218_));
 sky130_fd_sc_hd__or3_1 _13912_ (.A(_07536_),
    .B(_07527_),
    .C(_07528_),
    .X(_07538_));
 sky130_fd_sc_hd__or3_2 _13913_ (.A(_07518_),
    .B(_07538_),
    .C(_07501_),
    .X(_07539_));
 sky130_fd_sc_hd__nor2_1 _13914_ (.A(_07361_),
    .B(_07539_),
    .Y(_07540_));
 sky130_fd_sc_hd__or2_1 _13915_ (.A(\core.count_instr[40] ),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__buf_1 _13916_ (.A(_04388_),
    .X(_07542_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(_07540_),
    .B(\core.count_instr[40] ),
    .Y(_07543_));
 sky130_fd_sc_hd__and3_1 _13918_ (.A(_07541_),
    .B(_07542_),
    .C(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__buf_1 _13919_ (.A(_07544_),
    .X(_00219_));
 sky130_fd_sc_hd__or2_1 _13920_ (.A(\core.count_instr[41] ),
    .B(_07543_),
    .X(_07545_));
 sky130_fd_sc_hd__nand2_1 _13921_ (.A(_07543_),
    .B(\core.count_instr[41] ),
    .Y(_07546_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13922_ (.A(_04514_),
    .X(_07547_));
 sky130_fd_sc_hd__a21oi_1 _13923_ (.A1(_07545_),
    .A2(_07546_),
    .B1(_07547_),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _13924_ (.A(\core.count_instr[42] ),
    .Y(_07548_));
 sky130_fd_sc_hd__nand2_1 _13925_ (.A(\core.count_instr[41] ),
    .B(\core.count_instr[40] ),
    .Y(_07549_));
 sky130_fd_sc_hd__inv_2 _13926_ (.A(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__nand2_1 _13927_ (.A(_07540_),
    .B(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__nor2_1 _13928_ (.A(_07548_),
    .B(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__inv_2 _13929_ (.A(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__nand2_1 _13930_ (.A(_07551_),
    .B(_07548_),
    .Y(_07554_));
 sky130_fd_sc_hd__and3_1 _13931_ (.A(_07553_),
    .B(_07542_),
    .C(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__buf_1 _13932_ (.A(_07555_),
    .X(_00221_));
 sky130_fd_sc_hd__or2_1 _13933_ (.A(\core.count_instr[43] ),
    .B(_07553_),
    .X(_07556_));
 sky130_fd_sc_hd__nand2_1 _13934_ (.A(_07553_),
    .B(\core.count_instr[43] ),
    .Y(_07557_));
 sky130_fd_sc_hd__a21oi_1 _13935_ (.A1(_07556_),
    .A2(_07557_),
    .B1(_07547_),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _13936_ (.A(\core.count_instr[44] ),
    .Y(_07558_));
 sky130_fd_sc_hd__nor2_1 _13937_ (.A(_07518_),
    .B(_07538_),
    .Y(_07559_));
 sky130_fd_sc_hd__and3_1 _13938_ (.A(_07550_),
    .B(\core.count_instr[43] ),
    .C(\core.count_instr[42] ),
    .X(_07560_));
 sky130_fd_sc_hd__and4_1 _13939_ (.A(_07447_),
    .B(_07500_),
    .C(_07559_),
    .D(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__nand2_1 _13940_ (.A(_07561_),
    .B(_07414_),
    .Y(_07562_));
 sky130_fd_sc_hd__nor2_1 _13941_ (.A(_07558_),
    .B(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__inv_2 _13942_ (.A(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__nand2_1 _13943_ (.A(_07562_),
    .B(_07558_),
    .Y(_07565_));
 sky130_fd_sc_hd__and3_1 _13944_ (.A(_07564_),
    .B(_07542_),
    .C(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__clkbuf_1 _13945_ (.A(_07566_),
    .X(_00223_));
 sky130_fd_sc_hd__or2_1 _13946_ (.A(\core.count_instr[45] ),
    .B(_07564_),
    .X(_07567_));
 sky130_fd_sc_hd__nand2_1 _13947_ (.A(_07564_),
    .B(\core.count_instr[45] ),
    .Y(_07568_));
 sky130_fd_sc_hd__a21oi_1 _13948_ (.A1(_07567_),
    .A2(_07568_),
    .B1(_07547_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _13949_ (.A(\core.count_instr[45] ),
    .B(\core.count_instr[44] ),
    .Y(_07569_));
 sky130_fd_sc_hd__nor2_1 _13950_ (.A(_07569_),
    .B(_07562_),
    .Y(_07570_));
 sky130_fd_sc_hd__or2_2 _13951_ (.A(\core.count_instr[46] ),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__nand2_1 _13952_ (.A(_07570_),
    .B(\core.count_instr[46] ),
    .Y(_07572_));
 sky130_fd_sc_hd__and3_1 _13953_ (.A(_07571_),
    .B(_07542_),
    .C(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__buf_1 _13954_ (.A(_07573_),
    .X(_00225_));
 sky130_fd_sc_hd__or2_1 _13955_ (.A(\core.count_instr[47] ),
    .B(_07572_),
    .X(_07574_));
 sky130_fd_sc_hd__nand2_2 _13956_ (.A(_07572_),
    .B(\core.count_instr[47] ),
    .Y(_07575_));
 sky130_fd_sc_hd__a21oi_1 _13957_ (.A1(_07574_),
    .A2(_07575_),
    .B1(_07547_),
    .Y(_00226_));
 sky130_fd_sc_hd__and4_1 _13958_ (.A(\core.count_instr[47] ),
    .B(\core.count_instr[46] ),
    .C(\core.count_instr[45] ),
    .D(\core.count_instr[44] ),
    .X(_07576_));
 sky130_fd_sc_hd__and3_1 _13959_ (.A(_07559_),
    .B(_07560_),
    .C(_07576_),
    .X(_07577_));
 sky130_fd_sc_hd__and2_1 _13960_ (.A(_07415_),
    .B(_07431_),
    .X(_07578_));
 sky130_fd_sc_hd__and4_2 _13961_ (.A(_07399_),
    .B(_07577_),
    .C(_07500_),
    .D(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__nand2_4 _13962_ (.A(_07579_),
    .B(_07414_),
    .Y(_07580_));
 sky130_fd_sc_hd__inv_2 _13963_ (.A(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__or2_1 _13964_ (.A(\core.count_instr[48] ),
    .B(_07581_),
    .X(_07582_));
 sky130_fd_sc_hd__nand2_1 _13965_ (.A(_07581_),
    .B(\core.count_instr[48] ),
    .Y(_07583_));
 sky130_fd_sc_hd__and3_1 _13966_ (.A(_07582_),
    .B(_07542_),
    .C(_07583_),
    .X(_07584_));
 sky130_fd_sc_hd__clkbuf_1 _13967_ (.A(_07584_),
    .X(_00227_));
 sky130_fd_sc_hd__or2_1 _13968_ (.A(\core.count_instr[49] ),
    .B(_07583_),
    .X(_07585_));
 sky130_fd_sc_hd__nand2_1 _13969_ (.A(_07583_),
    .B(\core.count_instr[49] ),
    .Y(_07586_));
 sky130_fd_sc_hd__a21oi_1 _13970_ (.A1(_07585_),
    .A2(_07586_),
    .B1(_07547_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_2 _13971_ (.A(\core.count_instr[49] ),
    .B(\core.count_instr[48] ),
    .Y(_07587_));
 sky130_fd_sc_hd__nor2_2 _13972_ (.A(_07587_),
    .B(_07580_),
    .Y(_07588_));
 sky130_fd_sc_hd__or2_1 _13973_ (.A(\core.count_instr[50] ),
    .B(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(_07588_),
    .B(\core.count_instr[50] ),
    .Y(_07590_));
 sky130_fd_sc_hd__and3_1 _13975_ (.A(_07589_),
    .B(_07542_),
    .C(_07590_),
    .X(_07591_));
 sky130_fd_sc_hd__buf_1 _13976_ (.A(_07591_),
    .X(_00229_));
 sky130_fd_sc_hd__or2_1 _13977_ (.A(\core.count_instr[51] ),
    .B(_07590_),
    .X(_07592_));
 sky130_fd_sc_hd__nand2_1 _13978_ (.A(_07590_),
    .B(\core.count_instr[51] ),
    .Y(_07593_));
 sky130_fd_sc_hd__a21oi_1 _13979_ (.A1(_07592_),
    .A2(_07593_),
    .B1(_07547_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_2 _13980_ (.A(\core.count_instr[51] ),
    .B(\core.count_instr[50] ),
    .Y(_07594_));
 sky130_fd_sc_hd__nor2_2 _13981_ (.A(_07587_),
    .B(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__inv_2 _13982_ (.A(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__nor2_1 _13983_ (.A(_07596_),
    .B(_07580_),
    .Y(_07597_));
 sky130_fd_sc_hd__or2_1 _13984_ (.A(\core.count_instr[52] ),
    .B(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__nand2_1 _13985_ (.A(_07597_),
    .B(\core.count_instr[52] ),
    .Y(_07599_));
 sky130_fd_sc_hd__and3_1 _13986_ (.A(_07598_),
    .B(_04451_),
    .C(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__clkbuf_1 _13987_ (.A(_07600_),
    .X(_00231_));
 sky130_fd_sc_hd__and4_1 _13988_ (.A(_07579_),
    .B(\core.count_instr[52] ),
    .C(_07363_),
    .D(_07595_),
    .X(_07601_));
 sky130_fd_sc_hd__xor2_1 _13989_ (.A(\core.count_instr[53] ),
    .B(_07601_),
    .X(_07602_));
 sky130_fd_sc_hd__and2_1 _13990_ (.A(_07602_),
    .B(_06506_),
    .X(_07603_));
 sky130_fd_sc_hd__clkbuf_1 _13991_ (.A(_07603_),
    .X(_00232_));
 sky130_fd_sc_hd__nand2_1 _13992_ (.A(\core.count_instr[53] ),
    .B(\core.count_instr[52] ),
    .Y(_07604_));
 sky130_fd_sc_hd__nand3b_2 _13993_ (.A_N(_07604_),
    .B(_07579_),
    .C(_07595_),
    .Y(_07605_));
 sky130_fd_sc_hd__nor2_1 _13994_ (.A(_07379_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__or2_1 _13995_ (.A(\core.count_instr[54] ),
    .B(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__nand2_1 _13996_ (.A(_07606_),
    .B(\core.count_instr[54] ),
    .Y(_07608_));
 sky130_fd_sc_hd__and3_1 _13997_ (.A(_07607_),
    .B(_04451_),
    .C(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__buf_1 _13998_ (.A(_07609_),
    .X(_00233_));
 sky130_fd_sc_hd__or2_1 _13999_ (.A(\core.count_instr[55] ),
    .B(_07608_),
    .X(_07610_));
 sky130_fd_sc_hd__nand2_1 _14000_ (.A(_07608_),
    .B(\core.count_instr[55] ),
    .Y(_07611_));
 sky130_fd_sc_hd__buf_2 _14001_ (.A(_04514_),
    .X(_07612_));
 sky130_fd_sc_hd__a21oi_1 _14002_ (.A1(_07610_),
    .A2(_07611_),
    .B1(_07612_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _14003_ (.A(\core.count_instr[55] ),
    .B(\core.count_instr[54] ),
    .Y(_07613_));
 sky130_fd_sc_hd__nor3_1 _14004_ (.A(_07379_),
    .B(_07613_),
    .C(_07605_),
    .Y(_07614_));
 sky130_fd_sc_hd__a21oi_1 _14005_ (.A1(_07614_),
    .A2(\core.count_instr[56] ),
    .B1(_06326_),
    .Y(_07615_));
 sky130_fd_sc_hd__o21a_1 _14006_ (.A1(\core.count_instr[56] ),
    .A2(net105),
    .B1(_07615_),
    .X(_00235_));
 sky130_fd_sc_hd__a21bo_1 _14007_ (.A1(net105),
    .A2(\core.count_instr[56] ),
    .B1_N(\core.count_instr[57] ),
    .X(_07616_));
 sky130_fd_sc_hd__nand3b_1 _14008_ (.A_N(\core.count_instr[57] ),
    .B(net105),
    .C(\core.count_instr[56] ),
    .Y(_07617_));
 sky130_fd_sc_hd__a21oi_1 _14009_ (.A1(_07616_),
    .A2(_07617_),
    .B1(_07612_),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _14010_ (.A(\core.count_instr[58] ),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_1 _14011_ (.A(\core.count_instr[57] ),
    .B(\core.count_instr[56] ),
    .Y(_07619_));
 sky130_fd_sc_hd__or4_1 _14012_ (.A(_07379_),
    .B(_07613_),
    .C(_07619_),
    .D(_07605_),
    .X(_07620_));
 sky130_fd_sc_hd__o21ai_1 _14013_ (.A1(_07618_),
    .A2(_07620_),
    .B1(_06506_),
    .Y(_07621_));
 sky130_fd_sc_hd__a21oi_1 _14014_ (.A1(_07618_),
    .A2(_07620_),
    .B1(_07621_),
    .Y(_00237_));
 sky130_fd_sc_hd__or3_1 _14015_ (.A(_07604_),
    .B(_07613_),
    .C(_07596_),
    .X(_07622_));
 sky130_fd_sc_hd__and2b_2 _14016_ (.A_N(_07622_),
    .B(_07579_),
    .X(_07623_));
 sky130_fd_sc_hd__inv_2 _14017_ (.A(_07619_),
    .Y(_07624_));
 sky130_fd_sc_hd__and3_1 _14018_ (.A(_07623_),
    .B(\core.count_instr[58] ),
    .C(_07624_),
    .X(_07625_));
 sky130_fd_sc_hd__xor2_1 _14019_ (.A(\core.count_instr[59] ),
    .B(_07625_),
    .X(_07626_));
 sky130_fd_sc_hd__nand2_1 _14020_ (.A(_07626_),
    .B(_07375_),
    .Y(_07627_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14021_ (.A(_07379_),
    .X(_07628_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_07628_),
    .B(\core.count_instr[59] ),
    .Y(_07629_));
 sky130_fd_sc_hd__a21oi_1 _14023_ (.A1(_07627_),
    .A2(_07629_),
    .B1(_07612_),
    .Y(_00238_));
 sky130_fd_sc_hd__and3_1 _14024_ (.A(_07624_),
    .B(\core.count_instr[59] ),
    .C(\core.count_instr[58] ),
    .X(_07630_));
 sky130_fd_sc_hd__nand2_2 _14025_ (.A(_07623_),
    .B(_07630_),
    .Y(_07631_));
 sky130_fd_sc_hd__or2_1 _14026_ (.A(\core.count_instr[60] ),
    .B(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(_07631_),
    .B(\core.count_instr[60] ),
    .Y(_07633_));
 sky130_fd_sc_hd__a21o_1 _14028_ (.A1(_07632_),
    .A2(_07633_),
    .B1(_07628_),
    .X(_07634_));
 sky130_fd_sc_hd__nand2_1 _14029_ (.A(_07628_),
    .B(\core.count_instr[60] ),
    .Y(_07635_));
 sky130_fd_sc_hd__a21oi_1 _14030_ (.A1(_07634_),
    .A2(_07635_),
    .B1(_07612_),
    .Y(_00239_));
 sky130_fd_sc_hd__and3_1 _14031_ (.A(_07623_),
    .B(\core.count_instr[60] ),
    .C(_07630_),
    .X(_07636_));
 sky130_fd_sc_hd__xor2_1 _14032_ (.A(\core.count_instr[61] ),
    .B(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__nand2_1 _14033_ (.A(_07637_),
    .B(_07375_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _14034_ (.A(_07628_),
    .B(\core.count_instr[61] ),
    .Y(_07639_));
 sky130_fd_sc_hd__a21oi_1 _14035_ (.A1(_07638_),
    .A2(_07639_),
    .B1(_07612_),
    .Y(_00240_));
 sky130_fd_sc_hd__and4_1 _14036_ (.A(_07623_),
    .B(\core.count_instr[61] ),
    .C(\core.count_instr[60] ),
    .D(_07630_),
    .X(_07640_));
 sky130_fd_sc_hd__xor2_1 _14037_ (.A(\core.count_instr[62] ),
    .B(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__nand2_1 _14038_ (.A(_07641_),
    .B(_07375_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand2_1 _14039_ (.A(_07628_),
    .B(\core.count_instr[62] ),
    .Y(_07643_));
 sky130_fd_sc_hd__a21oi_1 _14040_ (.A1(_07642_),
    .A2(_07643_),
    .B1(_07612_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _14041_ (.A(_07640_),
    .B(\core.count_instr[62] ),
    .Y(_07644_));
 sky130_fd_sc_hd__nand2_1 _14042_ (.A(_07644_),
    .B(\core.count_instr[63] ),
    .Y(_07645_));
 sky130_fd_sc_hd__nand3b_1 _14043_ (.A_N(\core.count_instr[63] ),
    .B(_07640_),
    .C(\core.count_instr[62] ),
    .Y(_07646_));
 sky130_fd_sc_hd__nand2_1 _14044_ (.A(_07645_),
    .B(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__nand2_1 _14045_ (.A(_07647_),
    .B(_07375_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand2_1 _14046_ (.A(_07628_),
    .B(\core.count_instr[63] ),
    .Y(_07649_));
 sky130_fd_sc_hd__buf_2 _14047_ (.A(_04514_),
    .X(_07650_));
 sky130_fd_sc_hd__a21oi_1 _14048_ (.A1(_07648_),
    .A2(_07649_),
    .B1(_07650_),
    .Y(_00242_));
 sky130_fd_sc_hd__clkbuf_4 _14049_ (.A(_06321_),
    .X(_07651_));
 sky130_fd_sc_hd__buf_2 _14050_ (.A(_07651_),
    .X(_07652_));
 sky130_fd_sc_hd__or2_1 _14051_ (.A(_05011_),
    .B(\core.decoded_imm[0] ),
    .X(_07653_));
 sky130_fd_sc_hd__a21o_1 _14052_ (.A1(_05026_),
    .A2(_06235_),
    .B1(_04627_),
    .X(_07654_));
 sky130_fd_sc_hd__inv_2 _14053_ (.A(_06233_),
    .Y(_07655_));
 sky130_fd_sc_hd__buf_1 _14054_ (.A(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__buf_2 _14055_ (.A(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__inv_2 _14056_ (.A(_04481_),
    .Y(_07658_));
 sky130_fd_sc_hd__buf_2 _14057_ (.A(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__buf_2 _14058_ (.A(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__o21ai_2 _14059_ (.A1(_04730_),
    .A2(_07657_),
    .B1(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__a32o_1 _14060_ (.A1(_06225_),
    .A2(_06077_),
    .A3(_07653_),
    .B1(_07654_),
    .B2(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14061_ (.A(_06245_),
    .X(_07663_));
 sky130_fd_sc_hd__clkbuf_2 _14062_ (.A(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__clkbuf_2 _14063_ (.A(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__clkbuf_2 _14064_ (.A(_06275_),
    .X(_07666_));
 sky130_fd_sc_hd__clkbuf_2 _14065_ (.A(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__mux2_1 _14066_ (.A0(\core.cpuregs[6][0] ),
    .A1(\core.cpuregs[7][0] ),
    .S(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__clkbuf_2 _14067_ (.A(_07666_),
    .X(_07669_));
 sky130_fd_sc_hd__mux2_1 _14068_ (.A0(\core.cpuregs[4][0] ),
    .A1(\core.cpuregs[5][0] ),
    .S(_07669_),
    .X(_07670_));
 sky130_fd_sc_hd__clkbuf_2 _14069_ (.A(_06279_),
    .X(_07671_));
 sky130_fd_sc_hd__clkbuf_2 _14070_ (.A(_07671_),
    .X(_07672_));
 sky130_fd_sc_hd__buf_4 _14071_ (.A(_06253_),
    .X(_07673_));
 sky130_fd_sc_hd__a21o_1 _14072_ (.A1(_07670_),
    .A2(_07672_),
    .B1(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__a21oi_1 _14073_ (.A1(_07665_),
    .A2(_07668_),
    .B1(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__mux2_4 _14074_ (.A0(\core.cpuregs[0][0] ),
    .A1(\core.cpuregs[1][0] ),
    .S(_07669_),
    .X(_07676_));
 sky130_fd_sc_hd__nand2_1 _14075_ (.A(_07676_),
    .B(_07672_),
    .Y(_07677_));
 sky130_fd_sc_hd__mux2_4 _14076_ (.A0(\core.cpuregs[2][0] ),
    .A1(\core.cpuregs[3][0] ),
    .S(_07669_),
    .X(_07678_));
 sky130_fd_sc_hd__nand2_1 _14077_ (.A(_07678_),
    .B(_07665_),
    .Y(_07679_));
 sky130_fd_sc_hd__clkbuf_2 _14078_ (.A(_06254_),
    .X(_07680_));
 sky130_fd_sc_hd__a31o_1 _14079_ (.A1(_07677_),
    .A2(_07679_),
    .A3(_07680_),
    .B1(_00008_),
    .X(_07681_));
 sky130_fd_sc_hd__buf_6 _14080_ (.A(_00005_),
    .X(_07682_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14081_ (.A(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__clkbuf_2 _14082_ (.A(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__mux2_1 _14083_ (.A0(\core.cpuregs[14][0] ),
    .A1(\core.cpuregs[15][0] ),
    .S(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__mux2_1 _14084_ (.A0(\core.cpuregs[12][0] ),
    .A1(\core.cpuregs[13][0] ),
    .S(_07684_),
    .X(_07686_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14085_ (.A(_06278_),
    .X(_07687_));
 sky130_fd_sc_hd__clkbuf_2 _14086_ (.A(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__mux2_1 _14087_ (.A0(_07685_),
    .A1(_07686_),
    .S(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__mux2_1 _14088_ (.A0(\core.cpuregs[10][0] ),
    .A1(\core.cpuregs[11][0] ),
    .S(_07684_),
    .X(_07690_));
 sky130_fd_sc_hd__buf_6 _14089_ (.A(_07682_),
    .X(_07691_));
 sky130_fd_sc_hd__clkbuf_2 _14090_ (.A(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(\core.cpuregs[8][0] ),
    .A1(\core.cpuregs[9][0] ),
    .S(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__clkbuf_2 _14092_ (.A(_07687_),
    .X(_07694_));
 sky130_fd_sc_hd__mux2_1 _14093_ (.A0(_07690_),
    .A1(_07693_),
    .S(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__clkbuf_2 _14094_ (.A(_06253_),
    .X(_07696_));
 sky130_fd_sc_hd__mux2_1 _14095_ (.A0(_07689_),
    .A1(_07695_),
    .S(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__a2bb2o_1 _14096_ (.A1_N(_07675_),
    .A2_N(_07681_),
    .B1(_00008_),
    .B2(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__mux2_1 _14097_ (.A0(\core.cpuregs[28][0] ),
    .A1(\core.cpuregs[29][0] ),
    .S(_07667_),
    .X(_07699_));
 sky130_fd_sc_hd__mux2_1 _14098_ (.A0(\core.cpuregs[30][0] ),
    .A1(\core.cpuregs[31][0] ),
    .S(_07669_),
    .X(_07700_));
 sky130_fd_sc_hd__a21o_1 _14099_ (.A1(_07700_),
    .A2(_07665_),
    .B1(_07696_),
    .X(_07701_));
 sky130_fd_sc_hd__a21oi_1 _14100_ (.A1(_07672_),
    .A2(_07699_),
    .B1(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__mux2_1 _14101_ (.A0(\core.cpuregs[24][0] ),
    .A1(\core.cpuregs[25][0] ),
    .S(_07669_),
    .X(_07703_));
 sky130_fd_sc_hd__nand2_1 _14102_ (.A(_07703_),
    .B(_07672_),
    .Y(_07704_));
 sky130_fd_sc_hd__mux2_1 _14103_ (.A0(\core.cpuregs[26][0] ),
    .A1(\core.cpuregs[27][0] ),
    .S(_07669_),
    .X(_07705_));
 sky130_fd_sc_hd__nand2_1 _14104_ (.A(_07705_),
    .B(_07665_),
    .Y(_07706_));
 sky130_fd_sc_hd__a31o_1 _14105_ (.A1(_07704_),
    .A2(_07706_),
    .A3(_07680_),
    .B1(_06292_),
    .X(_07707_));
 sky130_fd_sc_hd__clkbuf_2 _14106_ (.A(_06292_),
    .X(_07708_));
 sky130_fd_sc_hd__mux2_4 _14107_ (.A0(\core.cpuregs[20][0] ),
    .A1(\core.cpuregs[21][0] ),
    .S(_07684_),
    .X(_07709_));
 sky130_fd_sc_hd__mux2_1 _14108_ (.A0(\core.cpuregs[22][0] ),
    .A1(\core.cpuregs[23][0] ),
    .S(_07692_),
    .X(_07710_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14109_ (.A(_06245_),
    .X(_07711_));
 sky130_fd_sc_hd__buf_4 _14110_ (.A(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__mux2_1 _14111_ (.A0(_07709_),
    .A1(_07710_),
    .S(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__mux2_1 _14112_ (.A0(\core.cpuregs[18][0] ),
    .A1(\core.cpuregs[19][0] ),
    .S(_07692_),
    .X(_07714_));
 sky130_fd_sc_hd__mux2_8 _14113_ (.A0(\core.cpuregs[16][0] ),
    .A1(\core.cpuregs[17][0] ),
    .S(_07692_),
    .X(_07715_));
 sky130_fd_sc_hd__mux2_1 _14114_ (.A0(_07714_),
    .A1(_07715_),
    .S(_07694_),
    .X(_07716_));
 sky130_fd_sc_hd__mux2_1 _14115_ (.A0(_07713_),
    .A1(_07716_),
    .S(_07696_),
    .X(_07717_));
 sky130_fd_sc_hd__a2bb2o_1 _14116_ (.A1_N(_07702_),
    .A2_N(_07707_),
    .B1(_07708_),
    .B2(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__buf_4 _14117_ (.A(_06268_),
    .X(_07719_));
 sky130_fd_sc_hd__clkbuf_4 _14118_ (.A(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__mux2_1 _14119_ (.A0(_07698_),
    .A1(_07718_),
    .S(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14120_ (.A(_06299_),
    .X(_07722_));
 sky130_fd_sc_hd__and3_1 _14121_ (.A(_07721_),
    .B(_06309_),
    .C(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__buf_1 _14122_ (.A(_06321_),
    .X(_07724_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14123_ (.A(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__o21ai_1 _14124_ (.A1(_07662_),
    .A2(_07723_),
    .B1(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__o21ai_2 _14125_ (.A1(_04693_),
    .A2(_07652_),
    .B1(_07726_),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _14126_ (.A(_06321_),
    .Y(_07727_));
 sky130_fd_sc_hd__clkbuf_2 _14127_ (.A(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__clkbuf_4 _14128_ (.A(_06301_),
    .X(_07729_));
 sky130_fd_sc_hd__nor2_1 _14129_ (.A(_07729_),
    .B(_05020_),
    .Y(_07730_));
 sky130_fd_sc_hd__buf_4 _14130_ (.A(_07666_),
    .X(_07731_));
 sky130_fd_sc_hd__mux2_1 _14131_ (.A0(\core.cpuregs[24][1] ),
    .A1(\core.cpuregs[25][1] ),
    .S(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(\core.cpuregs[26][1] ),
    .A1(\core.cpuregs[27][1] ),
    .S(_07731_),
    .X(_07733_));
 sky130_fd_sc_hd__mux2_1 _14133_ (.A0(_07732_),
    .A1(_07733_),
    .S(_07665_),
    .X(_07734_));
 sky130_fd_sc_hd__clkbuf_2 _14134_ (.A(_06254_),
    .X(_07735_));
 sky130_fd_sc_hd__nand2_1 _14135_ (.A(_07734_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__mux2_1 _14136_ (.A0(\core.cpuregs[28][1] ),
    .A1(\core.cpuregs[29][1] ),
    .S(_07731_),
    .X(_07737_));
 sky130_fd_sc_hd__mux2_1 _14137_ (.A0(\core.cpuregs[30][1] ),
    .A1(\core.cpuregs[31][1] ),
    .S(_07731_),
    .X(_07738_));
 sky130_fd_sc_hd__clkbuf_2 _14138_ (.A(_07663_),
    .X(_07739_));
 sky130_fd_sc_hd__mux2_4 _14139_ (.A0(_07737_),
    .A1(_07738_),
    .S(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__buf_2 _14140_ (.A(_06288_),
    .X(_07741_));
 sky130_fd_sc_hd__nand2_1 _14141_ (.A(_07740_),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14142_ (.A(_06275_),
    .X(_07743_));
 sky130_fd_sc_hd__clkbuf_2 _14143_ (.A(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__mux2_1 _14144_ (.A0(\core.cpuregs[12][1] ),
    .A1(\core.cpuregs[13][1] ),
    .S(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__clkbuf_2 _14145_ (.A(_07743_),
    .X(_07746_));
 sky130_fd_sc_hd__mux2_1 _14146_ (.A0(\core.cpuregs[14][1] ),
    .A1(\core.cpuregs[15][1] ),
    .S(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__mux2_1 _14147_ (.A0(_07745_),
    .A1(_07747_),
    .S(_07664_),
    .X(_07748_));
 sky130_fd_sc_hd__nand2_1 _14148_ (.A(_07748_),
    .B(_07741_),
    .Y(_07749_));
 sky130_fd_sc_hd__clkbuf_2 _14149_ (.A(_07743_),
    .X(_07750_));
 sky130_fd_sc_hd__mux2_1 _14150_ (.A0(\core.cpuregs[8][1] ),
    .A1(\core.cpuregs[9][1] ),
    .S(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__clkbuf_2 _14151_ (.A(_07743_),
    .X(_07752_));
 sky130_fd_sc_hd__mux2_1 _14152_ (.A0(\core.cpuregs[10][1] ),
    .A1(\core.cpuregs[11][1] ),
    .S(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__clkbuf_4 _14153_ (.A(_07663_),
    .X(_07754_));
 sky130_fd_sc_hd__mux2_1 _14154_ (.A0(_07751_),
    .A1(_07753_),
    .S(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__nand2_1 _14155_ (.A(_07755_),
    .B(_07735_),
    .Y(_07756_));
 sky130_fd_sc_hd__clkinv_4 _14156_ (.A(_06268_),
    .Y(_07757_));
 sky130_fd_sc_hd__and3_1 _14157_ (.A(_07749_),
    .B(_07756_),
    .C(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__a31o_1 _14158_ (.A1(_07719_),
    .A2(_07736_),
    .A3(_07742_),
    .B1(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__clkbuf_2 _14159_ (.A(_06298_),
    .X(_07760_));
 sky130_fd_sc_hd__a21oi_1 _14160_ (.A1(_07759_),
    .A2(_00008_),
    .B1(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__mux2_1 _14161_ (.A0(\core.cpuregs[16][1] ),
    .A1(\core.cpuregs[17][1] ),
    .S(_07667_),
    .X(_07762_));
 sky130_fd_sc_hd__mux2_4 _14162_ (.A0(\core.cpuregs[18][1] ),
    .A1(\core.cpuregs[19][1] ),
    .S(_07667_),
    .X(_07763_));
 sky130_fd_sc_hd__mux2_1 _14163_ (.A0(_07762_),
    .A1(_07763_),
    .S(_07665_),
    .X(_07764_));
 sky130_fd_sc_hd__nand2_1 _14164_ (.A(_07764_),
    .B(_07735_),
    .Y(_07765_));
 sky130_fd_sc_hd__mux2_1 _14165_ (.A0(\core.cpuregs[22][1] ),
    .A1(\core.cpuregs[23][1] ),
    .S(_07667_),
    .X(_07766_));
 sky130_fd_sc_hd__mux2_1 _14166_ (.A0(\core.cpuregs[20][1] ),
    .A1(\core.cpuregs[21][1] ),
    .S(_07667_),
    .X(_07767_));
 sky130_fd_sc_hd__mux2_2 _14167_ (.A0(_07766_),
    .A1(_07767_),
    .S(_07672_),
    .X(_07768_));
 sky130_fd_sc_hd__nand2_8 _14168_ (.A(_07768_),
    .B(_07741_),
    .Y(_07769_));
 sky130_fd_sc_hd__mux2_1 _14169_ (.A0(\core.cpuregs[6][1] ),
    .A1(\core.cpuregs[7][1] ),
    .S(_07731_),
    .X(_07770_));
 sky130_fd_sc_hd__mux2_1 _14170_ (.A0(\core.cpuregs[4][1] ),
    .A1(\core.cpuregs[5][1] ),
    .S(_07731_),
    .X(_07771_));
 sky130_fd_sc_hd__mux2_1 _14171_ (.A0(_07770_),
    .A1(_07771_),
    .S(_07672_),
    .X(_07772_));
 sky130_fd_sc_hd__clkbuf_2 _14172_ (.A(_07666_),
    .X(_07773_));
 sky130_fd_sc_hd__mux2_1 _14173_ (.A0(\core.cpuregs[0][1] ),
    .A1(\core.cpuregs[1][1] ),
    .S(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__mux2_1 _14174_ (.A0(\core.cpuregs[2][1] ),
    .A1(\core.cpuregs[3][1] ),
    .S(_07773_),
    .X(_07775_));
 sky130_fd_sc_hd__mux2_1 _14175_ (.A0(_07774_),
    .A1(_07775_),
    .S(_07739_),
    .X(_07776_));
 sky130_fd_sc_hd__and2_1 _14176_ (.A(_07776_),
    .B(_07735_),
    .X(_07777_));
 sky130_fd_sc_hd__a211oi_1 _14177_ (.A1(_07741_),
    .A2(_07772_),
    .B1(_07719_),
    .C1(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__a31o_1 _14178_ (.A1(_07719_),
    .A2(_07765_),
    .A3(_07769_),
    .B1(_07778_),
    .X(_07779_));
 sky130_fd_sc_hd__buf_4 _14179_ (.A(_07708_),
    .X(_07780_));
 sky130_fd_sc_hd__nand2_8 _14180_ (.A(_07779_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__a22o_1 _14181_ (.A1(\core.is_lui_auipc_jal ),
    .A2(_07730_),
    .B1(_07761_),
    .B2(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__clkbuf_2 _14182_ (.A(_06308_),
    .X(_07783_));
 sky130_fd_sc_hd__nand2_1 _14183_ (.A(_07782_),
    .B(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__nand2_1 _14184_ (.A(_06080_),
    .B(_06077_),
    .Y(_07785_));
 sky130_fd_sc_hd__clkbuf_2 _14185_ (.A(_07658_),
    .X(_07786_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14186_ (.A(_06234_),
    .X(_07787_));
 sky130_fd_sc_hd__nand2_1 _14187_ (.A(_07787_),
    .B(_04728_),
    .Y(_07788_));
 sky130_fd_sc_hd__a21oi_1 _14188_ (.A1(_07786_),
    .A2(_07788_),
    .B1(_06230_),
    .Y(_07789_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14189_ (.A(_07655_),
    .X(_07790_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14190_ (.A(_07655_),
    .X(_07791_));
 sky130_fd_sc_hd__nand2_1 _14191_ (.A(_07791_),
    .B(_04693_),
    .Y(_07792_));
 sky130_fd_sc_hd__o21ai_1 _14192_ (.A1(_04699_),
    .A2(_07790_),
    .B1(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand2_1 _14193_ (.A(_07793_),
    .B(_04626_),
    .Y(_07794_));
 sky130_fd_sc_hd__a32o_1 _14194_ (.A1(_04397_),
    .A2(_06082_),
    .A3(_07785_),
    .B1(_07789_),
    .B2(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__nor2_1 _14195_ (.A(_07795_),
    .B(_07727_),
    .Y(_07796_));
 sky130_fd_sc_hd__a22oi_2 _14196_ (.A1(_05049_),
    .A2(_07728_),
    .B1(_07784_),
    .B2(_07796_),
    .Y(_00244_));
 sky130_fd_sc_hd__or2_1 _14197_ (.A(_06090_),
    .B(_06083_),
    .X(_07797_));
 sky130_fd_sc_hd__nand2_1 _14198_ (.A(_06083_),
    .B(_06090_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_1 _14199_ (.A(_07655_),
    .B(_05032_),
    .Y(_07799_));
 sky130_fd_sc_hd__nand2_1 _14200_ (.A(_06234_),
    .B(_04700_),
    .Y(_07800_));
 sky130_fd_sc_hd__a21o_1 _14201_ (.A1(_07799_),
    .A2(_07800_),
    .B1(_07659_),
    .X(_07801_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14202_ (.A(_06233_),
    .X(_07802_));
 sky130_fd_sc_hd__nand2_1 _14203_ (.A(_07802_),
    .B(_04737_),
    .Y(_07803_));
 sky130_fd_sc_hd__a21oi_1 _14204_ (.A1(_07659_),
    .A2(_07803_),
    .B1(_04586_),
    .Y(_07804_));
 sky130_fd_sc_hd__a32o_1 _14205_ (.A1(_07797_),
    .A2(_04397_),
    .A3(_07798_),
    .B1(_07801_),
    .B2(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__or2_1 _14206_ (.A(_07805_),
    .B(_07727_),
    .X(_07806_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14207_ (.A(_06275_),
    .X(_07807_));
 sky130_fd_sc_hd__clkbuf_2 _14208_ (.A(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__mux2_1 _14209_ (.A0(\core.cpuregs[16][2] ),
    .A1(\core.cpuregs[17][2] ),
    .S(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__clkbuf_4 _14210_ (.A(_07807_),
    .X(_07810_));
 sky130_fd_sc_hd__mux2_1 _14211_ (.A0(\core.cpuregs[18][2] ),
    .A1(\core.cpuregs[19][2] ),
    .S(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__clkbuf_2 _14212_ (.A(_07663_),
    .X(_07812_));
 sky130_fd_sc_hd__mux2_1 _14213_ (.A0(_07809_),
    .A1(_07811_),
    .S(_07812_),
    .X(_07813_));
 sky130_fd_sc_hd__mux2_1 _14214_ (.A0(\core.cpuregs[22][2] ),
    .A1(\core.cpuregs[23][2] ),
    .S(_07810_),
    .X(_07814_));
 sky130_fd_sc_hd__mux2_1 _14215_ (.A0(\core.cpuregs[20][2] ),
    .A1(\core.cpuregs[21][2] ),
    .S(_07810_),
    .X(_07815_));
 sky130_fd_sc_hd__clkbuf_2 _14216_ (.A(_06279_),
    .X(_07816_));
 sky130_fd_sc_hd__mux2_1 _14217_ (.A0(_07814_),
    .A1(_07815_),
    .S(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__clkbuf_2 _14218_ (.A(_06288_),
    .X(_07818_));
 sky130_fd_sc_hd__mux2_1 _14219_ (.A0(_07813_),
    .A1(_07817_),
    .S(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__mux2_1 _14220_ (.A0(\core.cpuregs[24][2] ),
    .A1(\core.cpuregs[25][2] ),
    .S(_07808_),
    .X(_07820_));
 sky130_fd_sc_hd__mux2_1 _14221_ (.A0(\core.cpuregs[26][2] ),
    .A1(\core.cpuregs[27][2] ),
    .S(_07810_),
    .X(_07821_));
 sky130_fd_sc_hd__mux2_1 _14222_ (.A0(_07820_),
    .A1(_07821_),
    .S(_07812_),
    .X(_07822_));
 sky130_fd_sc_hd__mux2_1 _14223_ (.A0(\core.cpuregs[28][2] ),
    .A1(\core.cpuregs[29][2] ),
    .S(_07810_),
    .X(_07823_));
 sky130_fd_sc_hd__clkbuf_2 _14224_ (.A(_07807_),
    .X(_07824_));
 sky130_fd_sc_hd__mux2_1 _14225_ (.A0(\core.cpuregs[30][2] ),
    .A1(\core.cpuregs[31][2] ),
    .S(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__mux2_1 _14226_ (.A0(_07823_),
    .A1(_07825_),
    .S(_07812_),
    .X(_07826_));
 sky130_fd_sc_hd__clkbuf_4 _14227_ (.A(_00007_),
    .X(_07827_));
 sky130_fd_sc_hd__clkbuf_2 _14228_ (.A(_07827_),
    .X(_07828_));
 sky130_fd_sc_hd__mux2_1 _14229_ (.A0(_07822_),
    .A1(_07826_),
    .S(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__mux2_1 _14230_ (.A0(_07819_),
    .A1(_07829_),
    .S(_00008_),
    .X(_07830_));
 sky130_fd_sc_hd__mux2_1 _14231_ (.A0(\core.cpuregs[0][2] ),
    .A1(\core.cpuregs[1][2] ),
    .S(_07810_),
    .X(_07831_));
 sky130_fd_sc_hd__mux2_2 _14232_ (.A0(\core.cpuregs[2][2] ),
    .A1(\core.cpuregs[3][2] ),
    .S(_07824_),
    .X(_07832_));
 sky130_fd_sc_hd__mux2_1 _14233_ (.A0(_07831_),
    .A1(_07832_),
    .S(_07812_),
    .X(_07833_));
 sky130_fd_sc_hd__mux2_1 _14234_ (.A0(\core.cpuregs[6][2] ),
    .A1(\core.cpuregs[7][2] ),
    .S(_07824_),
    .X(_07834_));
 sky130_fd_sc_hd__clkbuf_2 _14235_ (.A(_07807_),
    .X(_07835_));
 sky130_fd_sc_hd__mux2_1 _14236_ (.A0(\core.cpuregs[4][2] ),
    .A1(\core.cpuregs[5][2] ),
    .S(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__mux2_1 _14237_ (.A0(_07834_),
    .A1(_07836_),
    .S(_07671_),
    .X(_07837_));
 sky130_fd_sc_hd__mux2_1 _14238_ (.A0(_07833_),
    .A1(_07837_),
    .S(_07828_),
    .X(_07838_));
 sky130_fd_sc_hd__mux2_1 _14239_ (.A0(\core.cpuregs[12][2] ),
    .A1(\core.cpuregs[13][2] ),
    .S(_07824_),
    .X(_07839_));
 sky130_fd_sc_hd__mux2_1 _14240_ (.A0(\core.cpuregs[14][2] ),
    .A1(\core.cpuregs[15][2] ),
    .S(_07824_),
    .X(_07840_));
 sky130_fd_sc_hd__clkbuf_2 _14241_ (.A(_07663_),
    .X(_07841_));
 sky130_fd_sc_hd__mux2_1 _14242_ (.A0(_07839_),
    .A1(_07840_),
    .S(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__mux2_1 _14243_ (.A0(\core.cpuregs[8][2] ),
    .A1(\core.cpuregs[9][2] ),
    .S(_07824_),
    .X(_07843_));
 sky130_fd_sc_hd__mux2_2 _14244_ (.A0(\core.cpuregs[10][2] ),
    .A1(\core.cpuregs[11][2] ),
    .S(_07835_),
    .X(_07844_));
 sky130_fd_sc_hd__mux2_1 _14245_ (.A0(_07843_),
    .A1(_07844_),
    .S(_07841_),
    .X(_07845_));
 sky130_fd_sc_hd__mux2_1 _14246_ (.A0(_07842_),
    .A1(_07845_),
    .S(_07680_),
    .X(_07846_));
 sky130_fd_sc_hd__mux2_1 _14247_ (.A0(_07838_),
    .A1(_07846_),
    .S(_00008_),
    .X(_07847_));
 sky130_fd_sc_hd__clkbuf_2 _14248_ (.A(_07757_),
    .X(_07848_));
 sky130_fd_sc_hd__mux2_1 _14249_ (.A0(_07830_),
    .A1(_07847_),
    .S(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__clkbuf_2 _14250_ (.A(_06299_),
    .X(_07850_));
 sky130_fd_sc_hd__nand2_1 _14251_ (.A(_07849_),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__buf_1 _14252_ (.A(_06304_),
    .X(_07852_));
 sky130_fd_sc_hd__or3_1 _14253_ (.A(_07729_),
    .B(_05053_),
    .C(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__inv_2 _14254_ (.A(_06308_),
    .Y(_07854_));
 sky130_fd_sc_hd__clkbuf_2 _14255_ (.A(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__a21oi_1 _14256_ (.A1(_07851_),
    .A2(_07853_),
    .B1(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__o22a_1 _14257_ (.A1(_04699_),
    .A2(_07652_),
    .B1(_07806_),
    .B2(_07856_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _14258_ (.A0(\core.cpuregs[24][3] ),
    .A1(\core.cpuregs[25][3] ),
    .S(_06276_),
    .X(_07857_));
 sky130_fd_sc_hd__clkbuf_4 _14259_ (.A(_06275_),
    .X(_07858_));
 sky130_fd_sc_hd__mux2_1 _14260_ (.A0(\core.cpuregs[26][3] ),
    .A1(\core.cpuregs[27][3] ),
    .S(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__buf_2 _14261_ (.A(_06245_),
    .X(_07860_));
 sky130_fd_sc_hd__mux2_1 _14262_ (.A0(_07857_),
    .A1(_07859_),
    .S(_07860_),
    .X(_07861_));
 sky130_fd_sc_hd__mux2_1 _14263_ (.A0(\core.cpuregs[28][3] ),
    .A1(\core.cpuregs[29][3] ),
    .S(_07858_),
    .X(_07862_));
 sky130_fd_sc_hd__mux2_1 _14264_ (.A0(\core.cpuregs[30][3] ),
    .A1(\core.cpuregs[31][3] ),
    .S(_07858_),
    .X(_07863_));
 sky130_fd_sc_hd__mux2_1 _14265_ (.A0(_07862_),
    .A1(_07863_),
    .S(_07860_),
    .X(_07864_));
 sky130_fd_sc_hd__mux2_1 _14266_ (.A0(_07861_),
    .A1(_07864_),
    .S(_06288_),
    .X(_07865_));
 sky130_fd_sc_hd__mux2_1 _14267_ (.A0(\core.cpuregs[16][3] ),
    .A1(\core.cpuregs[17][3] ),
    .S(_06276_),
    .X(_07866_));
 sky130_fd_sc_hd__mux2_1 _14268_ (.A0(\core.cpuregs[18][3] ),
    .A1(\core.cpuregs[19][3] ),
    .S(_07858_),
    .X(_07867_));
 sky130_fd_sc_hd__mux2_1 _14269_ (.A0(_07866_),
    .A1(_07867_),
    .S(_07860_),
    .X(_07868_));
 sky130_fd_sc_hd__mux2_1 _14270_ (.A0(\core.cpuregs[22][3] ),
    .A1(\core.cpuregs[23][3] ),
    .S(_07858_),
    .X(_07869_));
 sky130_fd_sc_hd__clkbuf_4 _14271_ (.A(_06275_),
    .X(_07870_));
 sky130_fd_sc_hd__mux2_1 _14272_ (.A0(\core.cpuregs[20][3] ),
    .A1(\core.cpuregs[21][3] ),
    .S(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__mux2_2 _14273_ (.A0(_07869_),
    .A1(_07871_),
    .S(_06279_),
    .X(_07872_));
 sky130_fd_sc_hd__mux2_1 _14274_ (.A0(_07868_),
    .A1(_07872_),
    .S(_06288_),
    .X(_07873_));
 sky130_fd_sc_hd__mux2_1 _14275_ (.A0(_07865_),
    .A1(_07873_),
    .S(_06292_),
    .X(_07874_));
 sky130_fd_sc_hd__mux2_1 _14276_ (.A0(\core.cpuregs[12][3] ),
    .A1(\core.cpuregs[13][3] ),
    .S(_07858_),
    .X(_07875_));
 sky130_fd_sc_hd__mux2_1 _14277_ (.A0(\core.cpuregs[14][3] ),
    .A1(\core.cpuregs[15][3] ),
    .S(_07870_),
    .X(_07876_));
 sky130_fd_sc_hd__mux2_1 _14278_ (.A0(_07875_),
    .A1(_07876_),
    .S(_07860_),
    .X(_07877_));
 sky130_fd_sc_hd__mux2_1 _14279_ (.A0(\core.cpuregs[8][3] ),
    .A1(\core.cpuregs[9][3] ),
    .S(_07870_),
    .X(_07878_));
 sky130_fd_sc_hd__mux2_1 _14280_ (.A0(\core.cpuregs[10][3] ),
    .A1(\core.cpuregs[11][3] ),
    .S(_07666_),
    .X(_07879_));
 sky130_fd_sc_hd__mux2_1 _14281_ (.A0(_07878_),
    .A1(_07879_),
    .S(_07860_),
    .X(_07880_));
 sky130_fd_sc_hd__mux2_1 _14282_ (.A0(_07877_),
    .A1(_07880_),
    .S(_06254_),
    .X(_07881_));
 sky130_fd_sc_hd__mux2_1 _14283_ (.A0(\core.cpuregs[0][3] ),
    .A1(\core.cpuregs[1][3] ),
    .S(_07870_),
    .X(_07882_));
 sky130_fd_sc_hd__mux2_1 _14284_ (.A0(\core.cpuregs[2][3] ),
    .A1(\core.cpuregs[3][3] ),
    .S(_07870_),
    .X(_07883_));
 sky130_fd_sc_hd__mux2_1 _14285_ (.A0(_07882_),
    .A1(_07883_),
    .S(_07860_),
    .X(_07884_));
 sky130_fd_sc_hd__mux2_1 _14286_ (.A0(\core.cpuregs[6][3] ),
    .A1(\core.cpuregs[7][3] ),
    .S(_07870_),
    .X(_07885_));
 sky130_fd_sc_hd__mux2_1 _14287_ (.A0(\core.cpuregs[4][3] ),
    .A1(\core.cpuregs[5][3] ),
    .S(_07666_),
    .X(_07886_));
 sky130_fd_sc_hd__mux2_1 _14288_ (.A0(_07885_),
    .A1(_07886_),
    .S(_06279_),
    .X(_07887_));
 sky130_fd_sc_hd__mux2_1 _14289_ (.A0(_07884_),
    .A1(_07887_),
    .S(_06288_),
    .X(_07888_));
 sky130_fd_sc_hd__mux2_2 _14290_ (.A0(_07881_),
    .A1(_07888_),
    .S(_06292_),
    .X(_07889_));
 sky130_fd_sc_hd__mux2_1 _14291_ (.A0(_07874_),
    .A1(_07889_),
    .S(_07757_),
    .X(_07890_));
 sky130_fd_sc_hd__nand2_1 _14292_ (.A(_07890_),
    .B(_06299_),
    .Y(_07891_));
 sky130_fd_sc_hd__buf_1 _14293_ (.A(_06304_),
    .X(_07892_));
 sky130_fd_sc_hd__or3b_1 _14294_ (.A(_06302_),
    .B(_07892_),
    .C_N(\core.reg_pc[3] ),
    .X(_07893_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14295_ (.A(_07854_),
    .X(_07894_));
 sky130_fd_sc_hd__a21o_1 _14296_ (.A1(_07891_),
    .A2(_07893_),
    .B1(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__a21o_1 _14297_ (.A1(_07798_),
    .A2(_06089_),
    .B1(_06086_),
    .X(_07896_));
 sky130_fd_sc_hd__nand2_1 _14298_ (.A(_07896_),
    .B(_04397_),
    .Y(_07897_));
 sky130_fd_sc_hd__a31o_1 _14299_ (.A1(_06086_),
    .A2(_06089_),
    .A3(_07798_),
    .B1(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__nand2_1 _14300_ (.A(_07655_),
    .B(_04683_),
    .Y(_07899_));
 sky130_fd_sc_hd__o21ai_1 _14301_ (.A1(_04723_),
    .A2(_07656_),
    .B1(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14302_ (.A(_06234_),
    .X(_07901_));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(_04481_),
    .X(_07902_));
 sky130_fd_sc_hd__a21oi_2 _14304_ (.A1(_07901_),
    .A2(_04734_),
    .B1(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__a211o_1 _14305_ (.A1(_07900_),
    .A2(_04626_),
    .B1(_04586_),
    .C1(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__and3_1 _14306_ (.A(_06321_),
    .B(_07898_),
    .C(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__a22oi_2 _14307_ (.A1(_04700_),
    .A2(_07727_),
    .B1(_07895_),
    .B2(_07905_),
    .Y(_00246_));
 sky130_fd_sc_hd__clkbuf_2 _14308_ (.A(_07807_),
    .X(_07906_));
 sky130_fd_sc_hd__mux2_1 _14309_ (.A0(\core.cpuregs[12][4] ),
    .A1(\core.cpuregs[13][4] ),
    .S(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14310_ (.A(_07682_),
    .X(_07908_));
 sky130_fd_sc_hd__clkbuf_4 _14311_ (.A(_07908_),
    .X(_07909_));
 sky130_fd_sc_hd__mux2_1 _14312_ (.A0(\core.cpuregs[14][4] ),
    .A1(\core.cpuregs[15][4] ),
    .S(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(_07907_),
    .A1(_07910_),
    .S(_07841_),
    .X(_07911_));
 sky130_fd_sc_hd__clkbuf_4 _14314_ (.A(_07908_),
    .X(_07912_));
 sky130_fd_sc_hd__mux2_1 _14315_ (.A0(\core.cpuregs[8][4] ),
    .A1(\core.cpuregs[9][4] ),
    .S(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__clkbuf_2 _14316_ (.A(_07908_),
    .X(_07914_));
 sky130_fd_sc_hd__mux2_1 _14317_ (.A0(\core.cpuregs[10][4] ),
    .A1(\core.cpuregs[11][4] ),
    .S(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__clkbuf_4 _14318_ (.A(_07711_),
    .X(_07916_));
 sky130_fd_sc_hd__mux2_1 _14319_ (.A0(_07913_),
    .A1(_07915_),
    .S(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__mux2_1 _14320_ (.A0(_07911_),
    .A1(_07917_),
    .S(_07680_),
    .X(_07918_));
 sky130_fd_sc_hd__clkbuf_4 _14321_ (.A(_07807_),
    .X(_07919_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(\core.cpuregs[24][4] ),
    .A1(\core.cpuregs[25][4] ),
    .S(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14323_ (.A(_07682_),
    .X(_07921_));
 sky130_fd_sc_hd__clkbuf_4 _14324_ (.A(_07921_),
    .X(_07922_));
 sky130_fd_sc_hd__mux2_1 _14325_ (.A0(\core.cpuregs[26][4] ),
    .A1(\core.cpuregs[27][4] ),
    .S(_07922_),
    .X(_07923_));
 sky130_fd_sc_hd__clkbuf_2 _14326_ (.A(_07711_),
    .X(_07924_));
 sky130_fd_sc_hd__mux2_1 _14327_ (.A0(_07920_),
    .A1(_07923_),
    .S(_07924_),
    .X(_07925_));
 sky130_fd_sc_hd__clkbuf_2 _14328_ (.A(_07908_),
    .X(_07926_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(\core.cpuregs[28][4] ),
    .A1(\core.cpuregs[29][4] ),
    .S(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__buf_4 _14330_ (.A(_07921_),
    .X(_07928_));
 sky130_fd_sc_hd__mux2_1 _14331_ (.A0(\core.cpuregs[30][4] ),
    .A1(\core.cpuregs[31][4] ),
    .S(_07928_),
    .X(_07929_));
 sky130_fd_sc_hd__clkbuf_2 _14332_ (.A(_07711_),
    .X(_07930_));
 sky130_fd_sc_hd__mux2_1 _14333_ (.A0(_07927_),
    .A1(_07929_),
    .S(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__mux2_1 _14334_ (.A0(_07925_),
    .A1(_07931_),
    .S(_07828_),
    .X(_07932_));
 sky130_fd_sc_hd__mux2_1 _14335_ (.A0(_07918_),
    .A1(_07932_),
    .S(_07719_),
    .X(_07933_));
 sky130_fd_sc_hd__clkbuf_4 _14336_ (.A(_07908_),
    .X(_07934_));
 sky130_fd_sc_hd__mux2_1 _14337_ (.A0(\core.cpuregs[0][4] ),
    .A1(\core.cpuregs[1][4] ),
    .S(_07934_),
    .X(_07935_));
 sky130_fd_sc_hd__clkbuf_2 _14338_ (.A(_07921_),
    .X(_07936_));
 sky130_fd_sc_hd__mux2_1 _14339_ (.A0(\core.cpuregs[2][4] ),
    .A1(\core.cpuregs[3][4] ),
    .S(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__clkbuf_4 _14340_ (.A(_07711_),
    .X(_07938_));
 sky130_fd_sc_hd__mux2_1 _14341_ (.A0(_07935_),
    .A1(_07937_),
    .S(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__clkbuf_4 _14342_ (.A(_07921_),
    .X(_07940_));
 sky130_fd_sc_hd__mux2_1 _14343_ (.A0(\core.cpuregs[6][4] ),
    .A1(\core.cpuregs[7][4] ),
    .S(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__clkbuf_2 _14344_ (.A(_07683_),
    .X(_07942_));
 sky130_fd_sc_hd__mux2_1 _14345_ (.A0(\core.cpuregs[4][4] ),
    .A1(\core.cpuregs[5][4] ),
    .S(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__mux2_1 _14346_ (.A0(_07941_),
    .A1(_07943_),
    .S(_07671_),
    .X(_07944_));
 sky130_fd_sc_hd__clkbuf_4 _14347_ (.A(_07827_),
    .X(_07945_));
 sky130_fd_sc_hd__mux2_1 _14348_ (.A0(_07939_),
    .A1(_07944_),
    .S(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__clkbuf_2 _14349_ (.A(_07921_),
    .X(_07947_));
 sky130_fd_sc_hd__mux2_1 _14350_ (.A0(\core.cpuregs[16][4] ),
    .A1(\core.cpuregs[17][4] ),
    .S(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__clkbuf_2 _14351_ (.A(_07683_),
    .X(_07949_));
 sky130_fd_sc_hd__mux2_1 _14352_ (.A0(\core.cpuregs[18][4] ),
    .A1(\core.cpuregs[19][4] ),
    .S(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__clkbuf_2 _14353_ (.A(_07711_),
    .X(_07951_));
 sky130_fd_sc_hd__mux2_1 _14354_ (.A0(_07948_),
    .A1(_07950_),
    .S(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__clkbuf_2 _14355_ (.A(_07683_),
    .X(_07953_));
 sky130_fd_sc_hd__mux2_1 _14356_ (.A0(\core.cpuregs[22][4] ),
    .A1(\core.cpuregs[23][4] ),
    .S(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__buf_2 _14357_ (.A(_07683_),
    .X(_07955_));
 sky130_fd_sc_hd__mux2_1 _14358_ (.A0(\core.cpuregs[20][4] ),
    .A1(\core.cpuregs[21][4] ),
    .S(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__clkbuf_2 _14359_ (.A(_07687_),
    .X(_07957_));
 sky130_fd_sc_hd__mux2_1 _14360_ (.A0(_07954_),
    .A1(_07956_),
    .S(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__clkbuf_4 _14361_ (.A(_07827_),
    .X(_07959_));
 sky130_fd_sc_hd__mux2_1 _14362_ (.A0(_07952_),
    .A1(_07958_),
    .S(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__buf_2 _14363_ (.A(_00009_),
    .X(_07961_));
 sky130_fd_sc_hd__mux2_1 _14364_ (.A0(_07946_),
    .A1(_07960_),
    .S(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__mux2_1 _14365_ (.A0(_07933_),
    .A1(_07962_),
    .S(_07780_),
    .X(_07963_));
 sky130_fd_sc_hd__buf_2 _14366_ (.A(\core.instr_lui ),
    .X(_07964_));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(\core.reg_pc[4] ),
    .Y(_07965_));
 sky130_fd_sc_hd__or3_2 _14368_ (.A(_07964_),
    .B(_07965_),
    .C(_07892_),
    .X(_07966_));
 sky130_fd_sc_hd__a21boi_2 _14369_ (.A1(_07963_),
    .A2(_07850_),
    .B1_N(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand2_1 _14370_ (.A(_07790_),
    .B(_04700_),
    .Y(_07968_));
 sky130_fd_sc_hd__nand2_1 _14371_ (.A(_07787_),
    .B(_04729_),
    .Y(_07969_));
 sky130_fd_sc_hd__clkbuf_2 _14372_ (.A(_07659_),
    .X(_07970_));
 sky130_fd_sc_hd__a21oi_2 _14373_ (.A1(_07968_),
    .A2(_07969_),
    .B1(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__nand2_1 _14374_ (.A(_07901_),
    .B(_04783_),
    .Y(_07972_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14375_ (.A(_07902_),
    .X(_07973_));
 sky130_fd_sc_hd__a21oi_2 _14376_ (.A1(_07792_),
    .A2(_07972_),
    .B1(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__nand2_1 _14377_ (.A(_06067_),
    .B(_06066_),
    .Y(_07975_));
 sky130_fd_sc_hd__nor2_1 _14378_ (.A(_07975_),
    .B(_06094_),
    .Y(_07976_));
 sky130_fd_sc_hd__a31o_1 _14379_ (.A1(_06091_),
    .A2(_06092_),
    .A3(_07975_),
    .B1(_04395_),
    .X(_07977_));
 sky130_fd_sc_hd__o32a_1 _14380_ (.A1(_04588_),
    .A2(_07971_),
    .A3(_07974_),
    .B1(_07976_),
    .B2(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__o21ai_2 _14381_ (.A1(_07855_),
    .A2(_07967_),
    .B1(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14382_ (.A(_07724_),
    .X(_07980_));
 sky130_fd_sc_hd__nand2_2 _14383_ (.A(_07979_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__o21ai_1 _14384_ (.A1(_04730_),
    .A2(_07652_),
    .B1(_07981_),
    .Y(_00247_));
 sky130_fd_sc_hd__mux2_1 _14385_ (.A0(\core.cpuregs[12][5] ),
    .A1(\core.cpuregs[13][5] ),
    .S(_07906_),
    .X(_07982_));
 sky130_fd_sc_hd__mux2_1 _14386_ (.A0(\core.cpuregs[14][5] ),
    .A1(\core.cpuregs[15][5] ),
    .S(_07909_),
    .X(_07983_));
 sky130_fd_sc_hd__buf_2 _14387_ (.A(_07663_),
    .X(_07984_));
 sky130_fd_sc_hd__mux2_1 _14388_ (.A0(_07982_),
    .A1(_07983_),
    .S(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__mux2_1 _14389_ (.A0(\core.cpuregs[8][5] ),
    .A1(\core.cpuregs[9][5] ),
    .S(_07912_),
    .X(_07986_));
 sky130_fd_sc_hd__mux2_1 _14390_ (.A0(\core.cpuregs[10][5] ),
    .A1(\core.cpuregs[11][5] ),
    .S(_07914_),
    .X(_07987_));
 sky130_fd_sc_hd__mux2_1 _14391_ (.A0(_07986_),
    .A1(_07987_),
    .S(_07916_),
    .X(_07988_));
 sky130_fd_sc_hd__mux2_1 _14392_ (.A0(_07985_),
    .A1(_07988_),
    .S(_07680_),
    .X(_07989_));
 sky130_fd_sc_hd__mux2_1 _14393_ (.A0(\core.cpuregs[24][5] ),
    .A1(\core.cpuregs[25][5] ),
    .S(_07912_),
    .X(_07990_));
 sky130_fd_sc_hd__clkbuf_4 _14394_ (.A(_07921_),
    .X(_07991_));
 sky130_fd_sc_hd__mux2_1 _14395_ (.A0(\core.cpuregs[26][5] ),
    .A1(\core.cpuregs[27][5] ),
    .S(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__mux2_1 _14396_ (.A0(_07990_),
    .A1(_07992_),
    .S(_07924_),
    .X(_07993_));
 sky130_fd_sc_hd__mux2_1 _14397_ (.A0(\core.cpuregs[28][5] ),
    .A1(\core.cpuregs[29][5] ),
    .S(_07926_),
    .X(_07994_));
 sky130_fd_sc_hd__mux2_1 _14398_ (.A0(\core.cpuregs[30][5] ),
    .A1(\core.cpuregs[31][5] ),
    .S(_07928_),
    .X(_07995_));
 sky130_fd_sc_hd__mux2_1 _14399_ (.A0(_07994_),
    .A1(_07995_),
    .S(_07930_),
    .X(_07996_));
 sky130_fd_sc_hd__mux2_1 _14400_ (.A0(_07993_),
    .A1(_07996_),
    .S(_07828_),
    .X(_07997_));
 sky130_fd_sc_hd__clkbuf_4 _14401_ (.A(_06268_),
    .X(_07998_));
 sky130_fd_sc_hd__mux2_1 _14402_ (.A0(_07989_),
    .A1(_07997_),
    .S(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__mux2_1 _14403_ (.A0(\core.cpuregs[0][5] ),
    .A1(\core.cpuregs[1][5] ),
    .S(_07934_),
    .X(_08000_));
 sky130_fd_sc_hd__mux2_1 _14404_ (.A0(\core.cpuregs[2][5] ),
    .A1(\core.cpuregs[3][5] ),
    .S(_07936_),
    .X(_08001_));
 sky130_fd_sc_hd__mux2_1 _14405_ (.A0(_08000_),
    .A1(_08001_),
    .S(_07938_),
    .X(_08002_));
 sky130_fd_sc_hd__mux2_1 _14406_ (.A0(\core.cpuregs[6][5] ),
    .A1(\core.cpuregs[7][5] ),
    .S(_07940_),
    .X(_08003_));
 sky130_fd_sc_hd__mux2_1 _14407_ (.A0(\core.cpuregs[4][5] ),
    .A1(\core.cpuregs[5][5] ),
    .S(_07942_),
    .X(_08004_));
 sky130_fd_sc_hd__mux2_1 _14408_ (.A0(_08003_),
    .A1(_08004_),
    .S(_07671_),
    .X(_08005_));
 sky130_fd_sc_hd__clkbuf_4 _14409_ (.A(_07827_),
    .X(_08006_));
 sky130_fd_sc_hd__mux2_1 _14410_ (.A0(_08002_),
    .A1(_08005_),
    .S(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__mux2_1 _14411_ (.A0(\core.cpuregs[16][5] ),
    .A1(\core.cpuregs[17][5] ),
    .S(_07947_),
    .X(_08008_));
 sky130_fd_sc_hd__clkbuf_4 _14412_ (.A(_07683_),
    .X(_08009_));
 sky130_fd_sc_hd__mux2_1 _14413_ (.A0(\core.cpuregs[18][5] ),
    .A1(\core.cpuregs[19][5] ),
    .S(_08009_),
    .X(_08010_));
 sky130_fd_sc_hd__mux2_1 _14414_ (.A0(_08008_),
    .A1(_08010_),
    .S(_07951_),
    .X(_08011_));
 sky130_fd_sc_hd__mux2_1 _14415_ (.A0(\core.cpuregs[22][5] ),
    .A1(\core.cpuregs[23][5] ),
    .S(_07953_),
    .X(_08012_));
 sky130_fd_sc_hd__mux2_1 _14416_ (.A0(\core.cpuregs[20][5] ),
    .A1(\core.cpuregs[21][5] ),
    .S(_07955_),
    .X(_08013_));
 sky130_fd_sc_hd__mux2_1 _14417_ (.A0(_08012_),
    .A1(_08013_),
    .S(_07957_),
    .X(_08014_));
 sky130_fd_sc_hd__mux2_1 _14418_ (.A0(_08011_),
    .A1(_08014_),
    .S(_07959_),
    .X(_08015_));
 sky130_fd_sc_hd__mux2_1 _14419_ (.A0(_08007_),
    .A1(_08015_),
    .S(_07961_),
    .X(_08016_));
 sky130_fd_sc_hd__mux2_1 _14420_ (.A0(_07999_),
    .A1(_08016_),
    .S(_07780_),
    .X(_08017_));
 sky130_fd_sc_hd__inv_2 _14421_ (.A(\core.reg_pc[5] ),
    .Y(_08018_));
 sky130_fd_sc_hd__or3_1 _14422_ (.A(_07964_),
    .B(_08018_),
    .C(_07892_),
    .X(_08019_));
 sky130_fd_sc_hd__a21boi_1 _14423_ (.A1(_08017_),
    .A2(_07850_),
    .B1_N(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand2_1 _14424_ (.A(_07791_),
    .B(_04730_),
    .Y(_08021_));
 sky130_fd_sc_hd__nand2_1 _14425_ (.A(_07787_),
    .B(_04738_),
    .Y(_08022_));
 sky130_fd_sc_hd__a21oi_1 _14426_ (.A1(_08021_),
    .A2(_08022_),
    .B1(_07970_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_1 _14427_ (.A(_07901_),
    .B(_04786_),
    .Y(_08024_));
 sky130_fd_sc_hd__a21oi_1 _14428_ (.A1(_07799_),
    .A2(_08024_),
    .B1(_07973_),
    .Y(_08025_));
 sky130_fd_sc_hd__o21ai_1 _14429_ (.A1(_07975_),
    .A2(_06094_),
    .B1(_06066_),
    .Y(_08026_));
 sky130_fd_sc_hd__or2_1 _14430_ (.A(_06065_),
    .B(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__nand2_1 _14431_ (.A(_08026_),
    .B(_06065_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _14432_ (.A(_08027_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__o32a_1 _14433_ (.A1(_04588_),
    .A2(_08023_),
    .A3(_08025_),
    .B1(_04984_),
    .B2(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__o21ai_1 _14434_ (.A1(_07855_),
    .A2(_08020_),
    .B1(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__nand2_1 _14435_ (.A(_08031_),
    .B(_07980_),
    .Y(_08032_));
 sky130_fd_sc_hd__o21ai_2 _14436_ (.A1(_04729_),
    .A2(_07652_),
    .B1(_08032_),
    .Y(_00248_));
 sky130_fd_sc_hd__buf_2 _14437_ (.A(_07651_),
    .X(_08033_));
 sky130_fd_sc_hd__mux2_1 _14438_ (.A0(\core.cpuregs[12][6] ),
    .A1(\core.cpuregs[13][6] ),
    .S(_07919_),
    .X(_08034_));
 sky130_fd_sc_hd__mux2_1 _14439_ (.A0(\core.cpuregs[14][6] ),
    .A1(\core.cpuregs[15][6] ),
    .S(_07909_),
    .X(_08035_));
 sky130_fd_sc_hd__mux2_1 _14440_ (.A0(_08034_),
    .A1(_08035_),
    .S(_07984_),
    .X(_08036_));
 sky130_fd_sc_hd__mux2_1 _14441_ (.A0(\core.cpuregs[8][6] ),
    .A1(\core.cpuregs[9][6] ),
    .S(_07912_),
    .X(_08037_));
 sky130_fd_sc_hd__mux2_1 _14442_ (.A0(\core.cpuregs[10][6] ),
    .A1(\core.cpuregs[11][6] ),
    .S(_07922_),
    .X(_08038_));
 sky130_fd_sc_hd__mux2_1 _14443_ (.A0(_08037_),
    .A1(_08038_),
    .S(_07916_),
    .X(_08039_));
 sky130_fd_sc_hd__mux2_1 _14444_ (.A0(_08036_),
    .A1(_08039_),
    .S(_07673_),
    .X(_08040_));
 sky130_fd_sc_hd__mux2_1 _14445_ (.A0(\core.cpuregs[24][6] ),
    .A1(\core.cpuregs[25][6] ),
    .S(_07912_),
    .X(_08041_));
 sky130_fd_sc_hd__mux2_2 _14446_ (.A0(\core.cpuregs[26][6] ),
    .A1(\core.cpuregs[27][6] ),
    .S(_07991_),
    .X(_08042_));
 sky130_fd_sc_hd__mux2_1 _14447_ (.A0(_08041_),
    .A1(_08042_),
    .S(_07924_),
    .X(_08043_));
 sky130_fd_sc_hd__mux2_1 _14448_ (.A0(\core.cpuregs[28][6] ),
    .A1(\core.cpuregs[29][6] ),
    .S(_07926_),
    .X(_08044_));
 sky130_fd_sc_hd__mux2_1 _14449_ (.A0(\core.cpuregs[30][6] ),
    .A1(\core.cpuregs[31][6] ),
    .S(_07928_),
    .X(_08045_));
 sky130_fd_sc_hd__mux2_1 _14450_ (.A0(_08044_),
    .A1(_08045_),
    .S(_07930_),
    .X(_08046_));
 sky130_fd_sc_hd__mux2_1 _14451_ (.A0(_08043_),
    .A1(_08046_),
    .S(_07945_),
    .X(_08047_));
 sky130_fd_sc_hd__mux2_1 _14452_ (.A0(_08040_),
    .A1(_08047_),
    .S(_07998_),
    .X(_08048_));
 sky130_fd_sc_hd__mux2_1 _14453_ (.A0(\core.cpuregs[0][6] ),
    .A1(\core.cpuregs[1][6] ),
    .S(_07934_),
    .X(_08049_));
 sky130_fd_sc_hd__mux2_1 _14454_ (.A0(\core.cpuregs[2][6] ),
    .A1(\core.cpuregs[3][6] ),
    .S(_07936_),
    .X(_08050_));
 sky130_fd_sc_hd__mux2_1 _14455_ (.A0(_08049_),
    .A1(_08050_),
    .S(_07938_),
    .X(_08051_));
 sky130_fd_sc_hd__mux2_1 _14456_ (.A0(\core.cpuregs[6][6] ),
    .A1(\core.cpuregs[7][6] ),
    .S(_07940_),
    .X(_08052_));
 sky130_fd_sc_hd__mux2_1 _14457_ (.A0(\core.cpuregs[4][6] ),
    .A1(\core.cpuregs[5][6] ),
    .S(_07942_),
    .X(_08053_));
 sky130_fd_sc_hd__mux2_1 _14458_ (.A0(_08052_),
    .A1(_08053_),
    .S(_07671_),
    .X(_08054_));
 sky130_fd_sc_hd__mux2_1 _14459_ (.A0(_08051_),
    .A1(_08054_),
    .S(_08006_),
    .X(_08055_));
 sky130_fd_sc_hd__mux2_1 _14460_ (.A0(\core.cpuregs[16][6] ),
    .A1(\core.cpuregs[17][6] ),
    .S(_07947_),
    .X(_08056_));
 sky130_fd_sc_hd__mux2_1 _14461_ (.A0(\core.cpuregs[18][6] ),
    .A1(\core.cpuregs[19][6] ),
    .S(_08009_),
    .X(_08057_));
 sky130_fd_sc_hd__mux2_1 _14462_ (.A0(_08056_),
    .A1(_08057_),
    .S(_07712_),
    .X(_08058_));
 sky130_fd_sc_hd__mux2_1 _14463_ (.A0(\core.cpuregs[22][6] ),
    .A1(\core.cpuregs[23][6] ),
    .S(_07949_),
    .X(_08059_));
 sky130_fd_sc_hd__mux2_1 _14464_ (.A0(\core.cpuregs[20][6] ),
    .A1(\core.cpuregs[21][6] ),
    .S(_07955_),
    .X(_08060_));
 sky130_fd_sc_hd__mux2_1 _14465_ (.A0(_08059_),
    .A1(_08060_),
    .S(_07688_),
    .X(_08061_));
 sky130_fd_sc_hd__mux2_1 _14466_ (.A0(_08058_),
    .A1(_08061_),
    .S(_07959_),
    .X(_08062_));
 sky130_fd_sc_hd__mux2_1 _14467_ (.A0(_08055_),
    .A1(_08062_),
    .S(_07961_),
    .X(_08063_));
 sky130_fd_sc_hd__mux2_1 _14468_ (.A0(_08048_),
    .A1(_08063_),
    .S(_07780_),
    .X(_08064_));
 sky130_fd_sc_hd__buf_1 _14469_ (.A(_06304_),
    .X(_08065_));
 sky130_fd_sc_hd__or3b_1 _14470_ (.A(_07964_),
    .B(_08065_),
    .C_N(_05122_),
    .X(_08066_));
 sky130_fd_sc_hd__a21boi_2 _14471_ (.A1(_08064_),
    .A2(_07850_),
    .B1_N(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__nand2_1 _14472_ (.A(_07791_),
    .B(_04729_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand2_1 _14473_ (.A(_07787_),
    .B(_04735_),
    .Y(_08069_));
 sky130_fd_sc_hd__a21oi_1 _14474_ (.A1(_08068_),
    .A2(_08069_),
    .B1(_07970_),
    .Y(_08070_));
 sky130_fd_sc_hd__nand2_1 _14475_ (.A(_07901_),
    .B(_04790_),
    .Y(_08071_));
 sky130_fd_sc_hd__a21oi_1 _14476_ (.A1(_07899_),
    .A2(_08071_),
    .B1(_07973_),
    .Y(_08072_));
 sky130_fd_sc_hd__a21o_1 _14477_ (.A1(_06093_),
    .A2(_06068_),
    .B1(_06096_),
    .X(_08073_));
 sky130_fd_sc_hd__or2_1 _14478_ (.A(_06074_),
    .B(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__nand2_1 _14479_ (.A(_08073_),
    .B(_06074_),
    .Y(_08075_));
 sky130_fd_sc_hd__nand2_4 _14480_ (.A(_08074_),
    .B(_08075_),
    .Y(_08076_));
 sky130_fd_sc_hd__o32a_1 _14481_ (.A1(_04588_),
    .A2(_08070_),
    .A3(_08072_),
    .B1(_04983_),
    .B2(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__o21ai_1 _14482_ (.A1(_07855_),
    .A2(_08067_),
    .B1(_08077_),
    .Y(_08078_));
 sky130_fd_sc_hd__nand2_1 _14483_ (.A(_08078_),
    .B(_07980_),
    .Y(_08079_));
 sky130_fd_sc_hd__o21ai_1 _14484_ (.A1(_04738_),
    .A2(_08033_),
    .B1(_08079_),
    .Y(_00249_));
 sky130_fd_sc_hd__mux2_1 _14485_ (.A0(\core.cpuregs[12][7] ),
    .A1(\core.cpuregs[13][7] ),
    .S(_07919_),
    .X(_08080_));
 sky130_fd_sc_hd__mux2_1 _14486_ (.A0(\core.cpuregs[14][7] ),
    .A1(\core.cpuregs[15][7] ),
    .S(_07909_),
    .X(_08081_));
 sky130_fd_sc_hd__mux2_1 _14487_ (.A0(_08080_),
    .A1(_08081_),
    .S(_07984_),
    .X(_08082_));
 sky130_fd_sc_hd__clkbuf_2 _14488_ (.A(_07908_),
    .X(_08083_));
 sky130_fd_sc_hd__mux2_1 _14489_ (.A0(\core.cpuregs[8][7] ),
    .A1(\core.cpuregs[9][7] ),
    .S(_08083_),
    .X(_08084_));
 sky130_fd_sc_hd__mux2_1 _14490_ (.A0(\core.cpuregs[10][7] ),
    .A1(\core.cpuregs[11][7] ),
    .S(_07922_),
    .X(_08085_));
 sky130_fd_sc_hd__mux2_1 _14491_ (.A0(_08084_),
    .A1(_08085_),
    .S(_07916_),
    .X(_08086_));
 sky130_fd_sc_hd__mux2_1 _14492_ (.A0(_08082_),
    .A1(_08086_),
    .S(_07673_),
    .X(_08087_));
 sky130_fd_sc_hd__mux2_1 _14493_ (.A0(\core.cpuregs[24][7] ),
    .A1(\core.cpuregs[25][7] ),
    .S(_07912_),
    .X(_08088_));
 sky130_fd_sc_hd__mux2_1 _14494_ (.A0(\core.cpuregs[26][7] ),
    .A1(\core.cpuregs[27][7] ),
    .S(_07991_),
    .X(_08089_));
 sky130_fd_sc_hd__mux2_1 _14495_ (.A0(_08088_),
    .A1(_08089_),
    .S(_07924_),
    .X(_08090_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(\core.cpuregs[28][7] ),
    .A1(\core.cpuregs[29][7] ),
    .S(_07914_),
    .X(_08091_));
 sky130_fd_sc_hd__mux2_1 _14497_ (.A0(\core.cpuregs[30][7] ),
    .A1(\core.cpuregs[31][7] ),
    .S(_07953_),
    .X(_08092_));
 sky130_fd_sc_hd__mux2_1 _14498_ (.A0(_08091_),
    .A1(_08092_),
    .S(_07951_),
    .X(_08093_));
 sky130_fd_sc_hd__mux2_1 _14499_ (.A0(_08090_),
    .A1(_08093_),
    .S(_07945_),
    .X(_08094_));
 sky130_fd_sc_hd__mux2_1 _14500_ (.A0(_08087_),
    .A1(_08094_),
    .S(_07998_),
    .X(_08095_));
 sky130_fd_sc_hd__mux2_1 _14501_ (.A0(\core.cpuregs[0][7] ),
    .A1(\core.cpuregs[1][7] ),
    .S(_07934_),
    .X(_08096_));
 sky130_fd_sc_hd__mux2_1 _14502_ (.A0(\core.cpuregs[2][7] ),
    .A1(\core.cpuregs[3][7] ),
    .S(_07936_),
    .X(_08097_));
 sky130_fd_sc_hd__mux2_1 _14503_ (.A0(_08096_),
    .A1(_08097_),
    .S(_07938_),
    .X(_08098_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(\core.cpuregs[6][7] ),
    .A1(\core.cpuregs[7][7] ),
    .S(_07940_),
    .X(_08099_));
 sky130_fd_sc_hd__mux2_1 _14505_ (.A0(\core.cpuregs[4][7] ),
    .A1(\core.cpuregs[5][7] ),
    .S(_07942_),
    .X(_08100_));
 sky130_fd_sc_hd__mux2_1 _14506_ (.A0(_08099_),
    .A1(_08100_),
    .S(_07957_),
    .X(_08101_));
 sky130_fd_sc_hd__mux2_1 _14507_ (.A0(_08098_),
    .A1(_08101_),
    .S(_08006_),
    .X(_08102_));
 sky130_fd_sc_hd__mux2_1 _14508_ (.A0(\core.cpuregs[16][7] ),
    .A1(\core.cpuregs[17][7] ),
    .S(_07947_),
    .X(_08103_));
 sky130_fd_sc_hd__mux2_1 _14509_ (.A0(\core.cpuregs[18][7] ),
    .A1(\core.cpuregs[19][7] ),
    .S(_08009_),
    .X(_08104_));
 sky130_fd_sc_hd__mux2_1 _14510_ (.A0(_08103_),
    .A1(_08104_),
    .S(_07712_),
    .X(_08105_));
 sky130_fd_sc_hd__mux2_2 _14511_ (.A0(\core.cpuregs[22][7] ),
    .A1(\core.cpuregs[23][7] ),
    .S(_07949_),
    .X(_08106_));
 sky130_fd_sc_hd__mux2_1 _14512_ (.A0(\core.cpuregs[20][7] ),
    .A1(\core.cpuregs[21][7] ),
    .S(_07955_),
    .X(_08107_));
 sky130_fd_sc_hd__mux2_1 _14513_ (.A0(_08106_),
    .A1(_08107_),
    .S(_07688_),
    .X(_08108_));
 sky130_fd_sc_hd__mux2_1 _14514_ (.A0(_08105_),
    .A1(_08108_),
    .S(_07959_),
    .X(_08109_));
 sky130_fd_sc_hd__mux2_1 _14515_ (.A0(_08102_),
    .A1(_08109_),
    .S(_07961_),
    .X(_08110_));
 sky130_fd_sc_hd__mux2_1 _14516_ (.A0(_08095_),
    .A1(_08110_),
    .S(_07780_),
    .X(_08111_));
 sky130_fd_sc_hd__inv_2 _14517_ (.A(\core.reg_pc[7] ),
    .Y(_08112_));
 sky130_fd_sc_hd__or3_1 _14518_ (.A(_07964_),
    .B(_08112_),
    .C(_07892_),
    .X(_08113_));
 sky130_fd_sc_hd__a21boi_1 _14519_ (.A1(_08111_),
    .A2(_07850_),
    .B1_N(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _14520_ (.A(_07791_),
    .B(_04738_),
    .Y(_08115_));
 sky130_fd_sc_hd__a21oi_1 _14521_ (.A1(_08115_),
    .A2(_07972_),
    .B1(_07970_),
    .Y(_08116_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14522_ (.A(_06234_),
    .X(_08117_));
 sky130_fd_sc_hd__nand2_1 _14523_ (.A(_08117_),
    .B(_04792_),
    .Y(_08118_));
 sky130_fd_sc_hd__a21oi_1 _14524_ (.A1(_07968_),
    .A2(_08118_),
    .B1(_07973_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand2_1 _14525_ (.A(_08075_),
    .B(_06073_),
    .Y(_08120_));
 sky130_fd_sc_hd__xnor2_1 _14526_ (.A(_06071_),
    .B(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__o32a_1 _14527_ (.A1(_06230_),
    .A2(_08116_),
    .A3(_08119_),
    .B1(_04983_),
    .B2(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__o21ai_1 _14528_ (.A1(_07855_),
    .A2(_08114_),
    .B1(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(_08123_),
    .B(_07980_),
    .Y(_08124_));
 sky130_fd_sc_hd__o21ai_1 _14530_ (.A1(_04735_),
    .A2(_08033_),
    .B1(_08124_),
    .Y(_00250_));
 sky130_fd_sc_hd__mux2_1 _14531_ (.A0(\core.cpuregs[12][8] ),
    .A1(\core.cpuregs[13][8] ),
    .S(_07919_),
    .X(_08125_));
 sky130_fd_sc_hd__mux2_1 _14532_ (.A0(\core.cpuregs[14][8] ),
    .A1(\core.cpuregs[15][8] ),
    .S(_07909_),
    .X(_08126_));
 sky130_fd_sc_hd__mux2_1 _14533_ (.A0(_08125_),
    .A1(_08126_),
    .S(_07984_),
    .X(_08127_));
 sky130_fd_sc_hd__mux2_1 _14534_ (.A0(\core.cpuregs[8][8] ),
    .A1(\core.cpuregs[9][8] ),
    .S(_08083_),
    .X(_08128_));
 sky130_fd_sc_hd__mux2_1 _14535_ (.A0(\core.cpuregs[10][8] ),
    .A1(\core.cpuregs[11][8] ),
    .S(_07922_),
    .X(_08129_));
 sky130_fd_sc_hd__mux2_1 _14536_ (.A0(_08128_),
    .A1(_08129_),
    .S(_07916_),
    .X(_08130_));
 sky130_fd_sc_hd__mux2_1 _14537_ (.A0(_08127_),
    .A1(_08130_),
    .S(_07673_),
    .X(_08131_));
 sky130_fd_sc_hd__mux2_1 _14538_ (.A0(\core.cpuregs[24][8] ),
    .A1(\core.cpuregs[25][8] ),
    .S(_08083_),
    .X(_08132_));
 sky130_fd_sc_hd__mux2_1 _14539_ (.A0(\core.cpuregs[26][8] ),
    .A1(\core.cpuregs[27][8] ),
    .S(_07991_),
    .X(_08133_));
 sky130_fd_sc_hd__mux2_2 _14540_ (.A0(_08132_),
    .A1(_08133_),
    .S(_07924_),
    .X(_08134_));
 sky130_fd_sc_hd__mux2_1 _14541_ (.A0(\core.cpuregs[28][8] ),
    .A1(\core.cpuregs[29][8] ),
    .S(_07914_),
    .X(_08135_));
 sky130_fd_sc_hd__mux2_2 _14542_ (.A0(\core.cpuregs[30][8] ),
    .A1(\core.cpuregs[31][8] ),
    .S(_07953_),
    .X(_08136_));
 sky130_fd_sc_hd__mux2_1 _14543_ (.A0(_08135_),
    .A1(_08136_),
    .S(_07951_),
    .X(_08137_));
 sky130_fd_sc_hd__mux2_1 _14544_ (.A0(_08134_),
    .A1(_08137_),
    .S(_07945_),
    .X(_08138_));
 sky130_fd_sc_hd__mux2_1 _14545_ (.A0(_08131_),
    .A1(_08138_),
    .S(_07998_),
    .X(_08139_));
 sky130_fd_sc_hd__mux2_1 _14546_ (.A0(\core.cpuregs[0][8] ),
    .A1(\core.cpuregs[1][8] ),
    .S(_07926_),
    .X(_08140_));
 sky130_fd_sc_hd__mux2_1 _14547_ (.A0(\core.cpuregs[2][8] ),
    .A1(\core.cpuregs[3][8] ),
    .S(_07928_),
    .X(_08141_));
 sky130_fd_sc_hd__mux2_4 _14548_ (.A0(_08140_),
    .A1(_08141_),
    .S(_07930_),
    .X(_08142_));
 sky130_fd_sc_hd__mux2_1 _14549_ (.A0(\core.cpuregs[6][8] ),
    .A1(\core.cpuregs[7][8] ),
    .S(_07940_),
    .X(_08143_));
 sky130_fd_sc_hd__mux2_1 _14550_ (.A0(\core.cpuregs[4][8] ),
    .A1(\core.cpuregs[5][8] ),
    .S(_07942_),
    .X(_08144_));
 sky130_fd_sc_hd__mux2_1 _14551_ (.A0(_08143_),
    .A1(_08144_),
    .S(_07957_),
    .X(_08145_));
 sky130_fd_sc_hd__mux2_1 _14552_ (.A0(_08142_),
    .A1(_08145_),
    .S(_08006_),
    .X(_08146_));
 sky130_fd_sc_hd__mux2_1 _14553_ (.A0(\core.cpuregs[16][8] ),
    .A1(\core.cpuregs[17][8] ),
    .S(_07947_),
    .X(_08147_));
 sky130_fd_sc_hd__mux2_1 _14554_ (.A0(\core.cpuregs[18][8] ),
    .A1(\core.cpuregs[19][8] ),
    .S(_08009_),
    .X(_08148_));
 sky130_fd_sc_hd__mux2_2 _14555_ (.A0(_08147_),
    .A1(_08148_),
    .S(_07712_),
    .X(_08149_));
 sky130_fd_sc_hd__mux2_2 _14556_ (.A0(\core.cpuregs[22][8] ),
    .A1(\core.cpuregs[23][8] ),
    .S(_07949_),
    .X(_08150_));
 sky130_fd_sc_hd__mux2_2 _14557_ (.A0(\core.cpuregs[20][8] ),
    .A1(\core.cpuregs[21][8] ),
    .S(_07955_),
    .X(_08151_));
 sky130_fd_sc_hd__mux2_1 _14558_ (.A0(_08150_),
    .A1(_08151_),
    .S(_07688_),
    .X(_08152_));
 sky130_fd_sc_hd__mux2_1 _14559_ (.A0(_08149_),
    .A1(_08152_),
    .S(_07959_),
    .X(_08153_));
 sky130_fd_sc_hd__mux2_1 _14560_ (.A0(_08146_),
    .A1(_08153_),
    .S(_07961_),
    .X(_08154_));
 sky130_fd_sc_hd__mux2_1 _14561_ (.A0(_08139_),
    .A1(_08154_),
    .S(_07780_),
    .X(_08155_));
 sky130_fd_sc_hd__inv_2 _14562_ (.A(\core.reg_pc[8] ),
    .Y(_08156_));
 sky130_fd_sc_hd__or3_1 _14563_ (.A(_07964_),
    .B(_08156_),
    .C(_07892_),
    .X(_08157_));
 sky130_fd_sc_hd__a21boi_1 _14564_ (.A1(_08155_),
    .A2(_07850_),
    .B1_N(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand2_1 _14565_ (.A(_07790_),
    .B(_04735_),
    .Y(_08159_));
 sky130_fd_sc_hd__a21oi_1 _14566_ (.A1(_08159_),
    .A2(_08024_),
    .B1(_07970_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_1 _14567_ (.A(_08117_),
    .B(_04796_),
    .Y(_08161_));
 sky130_fd_sc_hd__a21oi_1 _14568_ (.A1(_08021_),
    .A2(_08161_),
    .B1(_07973_),
    .Y(_08162_));
 sky130_fd_sc_hd__inv_2 _14569_ (.A(_06099_),
    .Y(_08163_));
 sky130_fd_sc_hd__nor2_1 _14570_ (.A(_06134_),
    .B(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__a21o_1 _14571_ (.A1(_08163_),
    .A2(_06134_),
    .B1(_04983_),
    .X(_08165_));
 sky130_fd_sc_hd__o32a_1 _14572_ (.A1(_06230_),
    .A2(_08160_),
    .A3(_08162_),
    .B1(_08164_),
    .B2(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__o21ai_1 _14573_ (.A1(_07855_),
    .A2(_08158_),
    .B1(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(_08167_),
    .B(_07980_),
    .Y(_08168_));
 sky130_fd_sc_hd__o21ai_2 _14575_ (.A1(_04783_),
    .A2(_08033_),
    .B1(_08168_),
    .Y(_00251_));
 sky130_fd_sc_hd__clkbuf_2 _14576_ (.A(_07854_),
    .X(_08169_));
 sky130_fd_sc_hd__mux2_1 _14577_ (.A0(\core.cpuregs[12][9] ),
    .A1(\core.cpuregs[13][9] ),
    .S(_07919_),
    .X(_08170_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\core.cpuregs[14][9] ),
    .A1(\core.cpuregs[15][9] ),
    .S(_07934_),
    .X(_08171_));
 sky130_fd_sc_hd__mux2_1 _14579_ (.A0(_08170_),
    .A1(_08171_),
    .S(_07984_),
    .X(_08172_));
 sky130_fd_sc_hd__mux2_1 _14580_ (.A0(\core.cpuregs[8][9] ),
    .A1(\core.cpuregs[9][9] ),
    .S(_08083_),
    .X(_08173_));
 sky130_fd_sc_hd__mux2_1 _14581_ (.A0(\core.cpuregs[10][9] ),
    .A1(\core.cpuregs[11][9] ),
    .S(_07922_),
    .X(_08174_));
 sky130_fd_sc_hd__mux2_1 _14582_ (.A0(_08173_),
    .A1(_08174_),
    .S(_07938_),
    .X(_08175_));
 sky130_fd_sc_hd__mux2_1 _14583_ (.A0(_08172_),
    .A1(_08175_),
    .S(_07673_),
    .X(_08176_));
 sky130_fd_sc_hd__mux2_1 _14584_ (.A0(\core.cpuregs[24][9] ),
    .A1(\core.cpuregs[25][9] ),
    .S(_08083_),
    .X(_08177_));
 sky130_fd_sc_hd__mux2_1 _14585_ (.A0(\core.cpuregs[26][9] ),
    .A1(\core.cpuregs[27][9] ),
    .S(_07991_),
    .X(_08178_));
 sky130_fd_sc_hd__mux2_1 _14586_ (.A0(_08177_),
    .A1(_08178_),
    .S(_07924_),
    .X(_08179_));
 sky130_fd_sc_hd__mux2_1 _14587_ (.A0(\core.cpuregs[28][9] ),
    .A1(\core.cpuregs[29][9] ),
    .S(_07914_),
    .X(_08180_));
 sky130_fd_sc_hd__mux2_1 _14588_ (.A0(\core.cpuregs[30][9] ),
    .A1(\core.cpuregs[31][9] ),
    .S(_07953_),
    .X(_08181_));
 sky130_fd_sc_hd__mux2_1 _14589_ (.A0(_08180_),
    .A1(_08181_),
    .S(_07951_),
    .X(_08182_));
 sky130_fd_sc_hd__mux2_1 _14590_ (.A0(_08179_),
    .A1(_08182_),
    .S(_07945_),
    .X(_08183_));
 sky130_fd_sc_hd__mux2_1 _14591_ (.A0(_08176_),
    .A1(_08183_),
    .S(_07998_),
    .X(_08184_));
 sky130_fd_sc_hd__mux2_1 _14592_ (.A0(\core.cpuregs[0][9] ),
    .A1(\core.cpuregs[1][9] ),
    .S(_07926_),
    .X(_08185_));
 sky130_fd_sc_hd__mux2_1 _14593_ (.A0(\core.cpuregs[2][9] ),
    .A1(\core.cpuregs[3][9] ),
    .S(_07928_),
    .X(_08186_));
 sky130_fd_sc_hd__mux2_2 _14594_ (.A0(_08185_),
    .A1(_08186_),
    .S(_07930_),
    .X(_08187_));
 sky130_fd_sc_hd__mux2_1 _14595_ (.A0(\core.cpuregs[6][9] ),
    .A1(\core.cpuregs[7][9] ),
    .S(_07936_),
    .X(_08188_));
 sky130_fd_sc_hd__mux2_1 _14596_ (.A0(\core.cpuregs[4][9] ),
    .A1(\core.cpuregs[5][9] ),
    .S(_07942_),
    .X(_08189_));
 sky130_fd_sc_hd__mux2_1 _14597_ (.A0(_08188_),
    .A1(_08189_),
    .S(_07957_),
    .X(_08190_));
 sky130_fd_sc_hd__mux2_1 _14598_ (.A0(_08187_),
    .A1(_08190_),
    .S(_08006_),
    .X(_08191_));
 sky130_fd_sc_hd__mux2_1 _14599_ (.A0(\core.cpuregs[16][9] ),
    .A1(\core.cpuregs[17][9] ),
    .S(_07947_),
    .X(_08192_));
 sky130_fd_sc_hd__mux2_1 _14600_ (.A0(\core.cpuregs[18][9] ),
    .A1(\core.cpuregs[19][9] ),
    .S(_08009_),
    .X(_08193_));
 sky130_fd_sc_hd__mux2_1 _14601_ (.A0(_08192_),
    .A1(_08193_),
    .S(_07712_),
    .X(_08194_));
 sky130_fd_sc_hd__mux2_1 _14602_ (.A0(\core.cpuregs[22][9] ),
    .A1(\core.cpuregs[23][9] ),
    .S(_07949_),
    .X(_08195_));
 sky130_fd_sc_hd__mux2_1 _14603_ (.A0(\core.cpuregs[20][9] ),
    .A1(\core.cpuregs[21][9] ),
    .S(_07684_),
    .X(_08196_));
 sky130_fd_sc_hd__mux2_1 _14604_ (.A0(_08195_),
    .A1(_08196_),
    .S(_07688_),
    .X(_08197_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(_08194_),
    .A1(_08197_),
    .S(_07959_),
    .X(_08198_));
 sky130_fd_sc_hd__mux2_1 _14606_ (.A0(_08191_),
    .A1(_08198_),
    .S(_07961_),
    .X(_08199_));
 sky130_fd_sc_hd__buf_2 _14607_ (.A(_06292_),
    .X(_08200_));
 sky130_fd_sc_hd__mux2_1 _14608_ (.A0(_08184_),
    .A1(_08199_),
    .S(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14609_ (.A(_06299_),
    .X(_08202_));
 sky130_fd_sc_hd__inv_2 _14610_ (.A(\core.reg_pc[9] ),
    .Y(_08203_));
 sky130_fd_sc_hd__or3_1 _14611_ (.A(_06301_),
    .B(_08203_),
    .C(_07892_),
    .X(_08204_));
 sky130_fd_sc_hd__a21boi_1 _14612_ (.A1(_08201_),
    .A2(_08202_),
    .B1_N(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nand2_1 _14613_ (.A(_07791_),
    .B(_04783_),
    .Y(_08206_));
 sky130_fd_sc_hd__a21oi_1 _14614_ (.A1(_08206_),
    .A2(_08071_),
    .B1(_07786_),
    .Y(_08207_));
 sky130_fd_sc_hd__nand2_1 _14615_ (.A(_07787_),
    .B(_04799_),
    .Y(_08208_));
 sky130_fd_sc_hd__a21oi_1 _14616_ (.A1(_08068_),
    .A2(_08208_),
    .B1(_07973_),
    .Y(_08209_));
 sky130_fd_sc_hd__o21a_1 _14617_ (.A1(_06134_),
    .A2(_08163_),
    .B1(_06133_),
    .X(_08210_));
 sky130_fd_sc_hd__nor2_1 _14618_ (.A(_06137_),
    .B(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(_08210_),
    .A2(_06137_),
    .B1(_04983_),
    .X(_08212_));
 sky130_fd_sc_hd__o32a_1 _14620_ (.A1(_06230_),
    .A2(_08207_),
    .A3(_08209_),
    .B1(_08211_),
    .B2(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__o21ai_1 _14621_ (.A1(_08169_),
    .A2(_08205_),
    .B1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14622_ (.A(_07724_),
    .X(_08215_));
 sky130_fd_sc_hd__nand2_1 _14623_ (.A(_08214_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__o21ai_2 _14624_ (.A1(_04786_),
    .A2(_08033_),
    .B1(_08216_),
    .Y(_00252_));
 sky130_fd_sc_hd__clkbuf_2 _14625_ (.A(_06239_),
    .X(_08217_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(\core.cpuregs[12][10] ),
    .A1(\core.cpuregs[13][10] ),
    .S(_08217_),
    .X(_08218_));
 sky130_fd_sc_hd__buf_4 _14627_ (.A(_06239_),
    .X(_08219_));
 sky130_fd_sc_hd__mux2_1 _14628_ (.A0(\core.cpuregs[14][10] ),
    .A1(\core.cpuregs[15][10] ),
    .S(_08219_),
    .X(_08220_));
 sky130_fd_sc_hd__clkbuf_2 _14629_ (.A(_06246_),
    .X(_08221_));
 sky130_fd_sc_hd__mux2_1 _14630_ (.A0(_08218_),
    .A1(_08220_),
    .S(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__mux2_1 _14631_ (.A0(\core.cpuregs[8][10] ),
    .A1(\core.cpuregs[9][10] ),
    .S(_08219_),
    .X(_08223_));
 sky130_fd_sc_hd__buf_4 _14632_ (.A(_06239_),
    .X(_08224_));
 sky130_fd_sc_hd__mux2_1 _14633_ (.A0(\core.cpuregs[10][10] ),
    .A1(\core.cpuregs[11][10] ),
    .S(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__clkbuf_2 _14634_ (.A(_06246_),
    .X(_08226_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(_08223_),
    .A1(_08225_),
    .S(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__mux2_1 _14636_ (.A0(_08222_),
    .A1(_08227_),
    .S(_06254_),
    .X(_08228_));
 sky130_fd_sc_hd__mux2_4 _14637_ (.A0(\core.cpuregs[24][10] ),
    .A1(\core.cpuregs[25][10] ),
    .S(_08219_),
    .X(_08229_));
 sky130_fd_sc_hd__clkbuf_2 _14638_ (.A(_06239_),
    .X(_08230_));
 sky130_fd_sc_hd__mux2_1 _14639_ (.A0(\core.cpuregs[26][10] ),
    .A1(\core.cpuregs[27][10] ),
    .S(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__mux2_1 _14640_ (.A0(_08229_),
    .A1(_08231_),
    .S(_08221_),
    .X(_08232_));
 sky130_fd_sc_hd__mux2_1 _14641_ (.A0(\core.cpuregs[28][10] ),
    .A1(\core.cpuregs[29][10] ),
    .S(_08224_),
    .X(_08233_));
 sky130_fd_sc_hd__buf_4 _14642_ (.A(_06239_),
    .X(_08234_));
 sky130_fd_sc_hd__mux2_1 _14643_ (.A0(\core.cpuregs[30][10] ),
    .A1(\core.cpuregs[31][10] ),
    .S(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__mux2_8 _14644_ (.A0(_08233_),
    .A1(_08235_),
    .S(_08226_),
    .X(_08236_));
 sky130_fd_sc_hd__buf_2 _14645_ (.A(_00007_),
    .X(_08237_));
 sky130_fd_sc_hd__clkbuf_2 _14646_ (.A(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__mux2_1 _14647_ (.A0(_08232_),
    .A1(_08236_),
    .S(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__clkbuf_2 _14648_ (.A(_00009_),
    .X(_08240_));
 sky130_fd_sc_hd__mux2_1 _14649_ (.A0(_08228_),
    .A1(_08239_),
    .S(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__mux2_4 _14650_ (.A0(\core.cpuregs[0][10] ),
    .A1(\core.cpuregs[1][10] ),
    .S(_08224_),
    .X(_08242_));
 sky130_fd_sc_hd__mux2_4 _14651_ (.A0(\core.cpuregs[2][10] ),
    .A1(\core.cpuregs[3][10] ),
    .S(_06240_),
    .X(_08243_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_08242_),
    .A1(_08243_),
    .S(_08226_),
    .X(_08244_));
 sky130_fd_sc_hd__mux2_1 _14653_ (.A0(\core.cpuregs[6][10] ),
    .A1(\core.cpuregs[7][10] ),
    .S(_08230_),
    .X(_08245_));
 sky130_fd_sc_hd__mux2_1 _14654_ (.A0(\core.cpuregs[4][10] ),
    .A1(\core.cpuregs[5][10] ),
    .S(_08234_),
    .X(_08246_));
 sky130_fd_sc_hd__clkbuf_2 _14655_ (.A(_06278_),
    .X(_08247_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(_08245_),
    .A1(_08246_),
    .S(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__clkbuf_2 _14657_ (.A(_08237_),
    .X(_08249_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(_08244_),
    .A1(_08248_),
    .S(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__mux2_8 _14659_ (.A0(\core.cpuregs[16][10] ),
    .A1(\core.cpuregs[17][10] ),
    .S(_08230_),
    .X(_08251_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(\core.cpuregs[18][10] ),
    .A1(\core.cpuregs[19][10] ),
    .S(_08234_),
    .X(_08252_));
 sky130_fd_sc_hd__clkbuf_2 _14661_ (.A(_06246_),
    .X(_08253_));
 sky130_fd_sc_hd__mux2_1 _14662_ (.A0(_08251_),
    .A1(_08252_),
    .S(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__mux2_1 _14663_ (.A0(\core.cpuregs[22][10] ),
    .A1(\core.cpuregs[23][10] ),
    .S(_08234_),
    .X(_08255_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(\core.cpuregs[20][10] ),
    .A1(\core.cpuregs[21][10] ),
    .S(_06260_),
    .X(_08256_));
 sky130_fd_sc_hd__clkbuf_2 _14665_ (.A(_06278_),
    .X(_08257_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(_08255_),
    .A1(_08256_),
    .S(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__mux2_4 _14667_ (.A0(_08254_),
    .A1(_08258_),
    .S(_08249_),
    .X(_08259_));
 sky130_fd_sc_hd__mux2_1 _14668_ (.A0(_08250_),
    .A1(_08259_),
    .S(_08240_),
    .X(_08260_));
 sky130_fd_sc_hd__mux2_1 _14669_ (.A0(_08241_),
    .A1(_08260_),
    .S(_06293_),
    .X(_08261_));
 sky130_fd_sc_hd__nand2_1 _14670_ (.A(_08261_),
    .B(_07722_),
    .Y(_08262_));
 sky130_fd_sc_hd__inv_2 _14671_ (.A(\core.reg_pc[10] ),
    .Y(_08263_));
 sky130_fd_sc_hd__or3_1 _14672_ (.A(_06302_),
    .B(_08263_),
    .C(_06305_),
    .X(_08264_));
 sky130_fd_sc_hd__a21o_1 _14673_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08169_),
    .X(_08265_));
 sky130_fd_sc_hd__a21bo_1 _14674_ (.A1(_06099_),
    .A2(_06138_),
    .B1_N(_06142_),
    .X(_08266_));
 sky130_fd_sc_hd__or2_1 _14675_ (.A(_06124_),
    .B(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__nand2_1 _14676_ (.A(_08266_),
    .B(_06124_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand3_1 _14677_ (.A(_08267_),
    .B(_06226_),
    .C(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14678_ (.A(_07656_),
    .X(_08270_));
 sky130_fd_sc_hd__nand2_1 _14679_ (.A(_08270_),
    .B(_04786_),
    .Y(_08271_));
 sky130_fd_sc_hd__clkbuf_2 _14680_ (.A(_07659_),
    .X(_08272_));
 sky130_fd_sc_hd__a21oi_2 _14681_ (.A1(_08271_),
    .A2(_08118_),
    .B1(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand2_1 _14682_ (.A(_08117_),
    .B(_04804_),
    .Y(_08274_));
 sky130_fd_sc_hd__a21oi_2 _14683_ (.A1(_08115_),
    .A2(_08274_),
    .B1(_04589_),
    .Y(_08275_));
 sky130_fd_sc_hd__o31a_1 _14684_ (.A1(_05319_),
    .A2(_08273_),
    .A3(_08275_),
    .B1(_07651_),
    .X(_08276_));
 sky130_fd_sc_hd__nand3_2 _14685_ (.A(_08265_),
    .B(_08269_),
    .C(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_2 _14686_ (.A(_07728_),
    .B(_04790_),
    .Y(_08278_));
 sky130_fd_sc_hd__nand2_8 _14687_ (.A(_08277_),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__inv_2 _14688_ (.A(_08279_),
    .Y(_00253_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14689_ (.A(_07682_),
    .X(_08280_));
 sky130_fd_sc_hd__buf_2 _14690_ (.A(_08280_),
    .X(_08281_));
 sky130_fd_sc_hd__mux2_1 _14691_ (.A0(\core.cpuregs[12][11] ),
    .A1(\core.cpuregs[13][11] ),
    .S(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__clkbuf_2 _14692_ (.A(_08280_),
    .X(_08283_));
 sky130_fd_sc_hd__mux2_1 _14693_ (.A0(\core.cpuregs[14][11] ),
    .A1(\core.cpuregs[15][11] ),
    .S(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14694_ (.A(_06245_),
    .X(_08285_));
 sky130_fd_sc_hd__clkbuf_4 _14695_ (.A(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__mux2_1 _14696_ (.A0(_08282_),
    .A1(_08284_),
    .S(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__clkbuf_2 _14697_ (.A(_08280_),
    .X(_08288_));
 sky130_fd_sc_hd__mux2_1 _14698_ (.A0(\core.cpuregs[8][11] ),
    .A1(\core.cpuregs[9][11] ),
    .S(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14699_ (.A(_06238_),
    .X(_08290_));
 sky130_fd_sc_hd__clkbuf_2 _14700_ (.A(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(\core.cpuregs[10][11] ),
    .A1(\core.cpuregs[11][11] ),
    .S(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14702_ (.A(_06245_),
    .X(_08293_));
 sky130_fd_sc_hd__clkbuf_4 _14703_ (.A(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__mux2_1 _14704_ (.A0(_08289_),
    .A1(_08292_),
    .S(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__clkbuf_2 _14705_ (.A(_06253_),
    .X(_08296_));
 sky130_fd_sc_hd__mux2_1 _14706_ (.A0(_08287_),
    .A1(_08295_),
    .S(_08296_),
    .X(_08297_));
 sky130_fd_sc_hd__clkbuf_2 _14707_ (.A(_08280_),
    .X(_08298_));
 sky130_fd_sc_hd__mux2_8 _14708_ (.A0(\core.cpuregs[24][11] ),
    .A1(\core.cpuregs[25][11] ),
    .S(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__clkbuf_2 _14709_ (.A(_08290_),
    .X(_08300_));
 sky130_fd_sc_hd__mux2_1 _14710_ (.A0(\core.cpuregs[26][11] ),
    .A1(\core.cpuregs[27][11] ),
    .S(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__clkbuf_2 _14711_ (.A(_08293_),
    .X(_08302_));
 sky130_fd_sc_hd__mux2_1 _14712_ (.A0(_08299_),
    .A1(_08301_),
    .S(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__clkbuf_2 _14713_ (.A(_08290_),
    .X(_08304_));
 sky130_fd_sc_hd__mux2_1 _14714_ (.A0(\core.cpuregs[28][11] ),
    .A1(\core.cpuregs[29][11] ),
    .S(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14715_ (.A(_06238_),
    .X(_08306_));
 sky130_fd_sc_hd__buf_4 _14716_ (.A(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(\core.cpuregs[30][11] ),
    .A1(\core.cpuregs[31][11] ),
    .S(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__clkbuf_2 _14718_ (.A(_08293_),
    .X(_08309_));
 sky130_fd_sc_hd__mux2_1 _14719_ (.A0(_08305_),
    .A1(_08308_),
    .S(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__buf_2 _14720_ (.A(_08237_),
    .X(_08311_));
 sky130_fd_sc_hd__mux2_1 _14721_ (.A0(_08303_),
    .A1(_08310_),
    .S(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__buf_2 _14722_ (.A(_00009_),
    .X(_08313_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(_08297_),
    .A1(_08312_),
    .S(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__clkbuf_4 _14724_ (.A(_08290_),
    .X(_08315_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(\core.cpuregs[0][11] ),
    .A1(\core.cpuregs[1][11] ),
    .S(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__clkbuf_4 _14726_ (.A(_08306_),
    .X(_08317_));
 sky130_fd_sc_hd__mux2_1 _14727_ (.A0(\core.cpuregs[2][11] ),
    .A1(\core.cpuregs[3][11] ),
    .S(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__clkbuf_4 _14728_ (.A(_08293_),
    .X(_08319_));
 sky130_fd_sc_hd__mux2_1 _14729_ (.A0(_08316_),
    .A1(_08318_),
    .S(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__clkbuf_4 _14730_ (.A(_08306_),
    .X(_08321_));
 sky130_fd_sc_hd__mux2_1 _14731_ (.A0(\core.cpuregs[6][11] ),
    .A1(\core.cpuregs[7][11] ),
    .S(_08321_),
    .X(_08322_));
 sky130_fd_sc_hd__clkbuf_2 _14732_ (.A(_08306_),
    .X(_08323_));
 sky130_fd_sc_hd__mux2_1 _14733_ (.A0(\core.cpuregs[4][11] ),
    .A1(\core.cpuregs[5][11] ),
    .S(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__clkbuf_2 _14734_ (.A(_07687_),
    .X(_08325_));
 sky130_fd_sc_hd__mux2_1 _14735_ (.A0(_08322_),
    .A1(_08324_),
    .S(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__clkbuf_2 _14736_ (.A(_08237_),
    .X(_08327_));
 sky130_fd_sc_hd__mux2_1 _14737_ (.A0(_08320_),
    .A1(_08326_),
    .S(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__clkbuf_2 _14738_ (.A(_08290_),
    .X(_08329_));
 sky130_fd_sc_hd__mux2_1 _14739_ (.A0(\core.cpuregs[16][11] ),
    .A1(\core.cpuregs[17][11] ),
    .S(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__mux2_1 _14740_ (.A0(\core.cpuregs[18][11] ),
    .A1(\core.cpuregs[19][11] ),
    .S(_08323_),
    .X(_08331_));
 sky130_fd_sc_hd__clkbuf_2 _14741_ (.A(_08293_),
    .X(_08332_));
 sky130_fd_sc_hd__mux2_1 _14742_ (.A0(_08330_),
    .A1(_08331_),
    .S(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__clkbuf_2 _14743_ (.A(_08306_),
    .X(_08334_));
 sky130_fd_sc_hd__mux2_1 _14744_ (.A0(\core.cpuregs[22][11] ),
    .A1(\core.cpuregs[23][11] ),
    .S(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14745_ (.A(_06238_),
    .X(_08336_));
 sky130_fd_sc_hd__clkbuf_2 _14746_ (.A(_08336_),
    .X(_08337_));
 sky130_fd_sc_hd__mux2_1 _14747_ (.A0(\core.cpuregs[20][11] ),
    .A1(\core.cpuregs[21][11] ),
    .S(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__clkbuf_2 _14748_ (.A(_07687_),
    .X(_08339_));
 sky130_fd_sc_hd__mux2_1 _14749_ (.A0(_08335_),
    .A1(_08338_),
    .S(_08339_),
    .X(_08340_));
 sky130_fd_sc_hd__clkbuf_2 _14750_ (.A(_08237_),
    .X(_08341_));
 sky130_fd_sc_hd__mux2_1 _14751_ (.A0(_08333_),
    .A1(_08340_),
    .S(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__clkbuf_2 _14752_ (.A(_00009_),
    .X(_08343_));
 sky130_fd_sc_hd__mux2_1 _14753_ (.A0(_08328_),
    .A1(_08342_),
    .S(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__mux2_1 _14754_ (.A0(_08314_),
    .A1(_08344_),
    .S(_08200_),
    .X(_08345_));
 sky130_fd_sc_hd__nand2_2 _14755_ (.A(_08345_),
    .B(_08202_),
    .Y(_08346_));
 sky130_fd_sc_hd__clkbuf_4 _14756_ (.A(_06301_),
    .X(_08347_));
 sky130_fd_sc_hd__inv_2 _14757_ (.A(\core.reg_pc[11] ),
    .Y(_08348_));
 sky130_fd_sc_hd__or3_1 _14758_ (.A(_08347_),
    .B(_08348_),
    .C(_07852_),
    .X(_08349_));
 sky130_fd_sc_hd__nand2_1 _14759_ (.A(_08346_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__nand2_1 _14760_ (.A(_08350_),
    .B(_07783_),
    .Y(_08351_));
 sky130_fd_sc_hd__a21oi_1 _14761_ (.A1(_08268_),
    .A2(_06122_),
    .B1(_06141_),
    .Y(_08352_));
 sky130_fd_sc_hd__a31o_1 _14762_ (.A1(_08268_),
    .A2(_06122_),
    .A3(_06141_),
    .B1(_04395_),
    .X(_08353_));
 sky130_fd_sc_hd__or2_1 _14763_ (.A(_08352_),
    .B(_08353_),
    .X(_08354_));
 sky130_fd_sc_hd__nand2_1 _14764_ (.A(_07657_),
    .B(_04790_),
    .Y(_08355_));
 sky130_fd_sc_hd__buf_1 _14765_ (.A(_07902_),
    .X(_08356_));
 sky130_fd_sc_hd__and3_1 _14766_ (.A(_08355_),
    .B(_08356_),
    .C(_08161_),
    .X(_08357_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14767_ (.A(_07802_),
    .X(_08358_));
 sky130_fd_sc_hd__nand2_1 _14768_ (.A(_08358_),
    .B(_04806_),
    .Y(_08359_));
 sky130_fd_sc_hd__and3_1 _14769_ (.A(_07660_),
    .B(_08159_),
    .C(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__o21ai_1 _14770_ (.A1(_08357_),
    .A2(_08360_),
    .B1(_04634_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand3_1 _14771_ (.A(_08351_),
    .B(_08354_),
    .C(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__nand2_1 _14772_ (.A(_08362_),
    .B(_08215_),
    .Y(_08363_));
 sky130_fd_sc_hd__o21ai_1 _14773_ (.A1(_04792_),
    .A2(_08033_),
    .B1(_08363_),
    .Y(_00254_));
 sky130_fd_sc_hd__mux2_1 _14774_ (.A0(\core.cpuregs[12][12] ),
    .A1(\core.cpuregs[13][12] ),
    .S(_08217_),
    .X(_08364_));
 sky130_fd_sc_hd__mux2_1 _14775_ (.A0(\core.cpuregs[14][12] ),
    .A1(\core.cpuregs[15][12] ),
    .S(_08219_),
    .X(_08365_));
 sky130_fd_sc_hd__mux2_1 _14776_ (.A0(_08364_),
    .A1(_08365_),
    .S(_08221_),
    .X(_08366_));
 sky130_fd_sc_hd__mux2_1 _14777_ (.A0(\core.cpuregs[8][12] ),
    .A1(\core.cpuregs[9][12] ),
    .S(_08219_),
    .X(_08367_));
 sky130_fd_sc_hd__mux2_1 _14778_ (.A0(\core.cpuregs[10][12] ),
    .A1(\core.cpuregs[11][12] ),
    .S(_08224_),
    .X(_08368_));
 sky130_fd_sc_hd__mux2_1 _14779_ (.A0(_08367_),
    .A1(_08368_),
    .S(_08226_),
    .X(_08369_));
 sky130_fd_sc_hd__mux2_1 _14780_ (.A0(_08366_),
    .A1(_08369_),
    .S(_06254_),
    .X(_08370_));
 sky130_fd_sc_hd__mux2_1 _14781_ (.A0(\core.cpuregs[24][12] ),
    .A1(\core.cpuregs[25][12] ),
    .S(_08219_),
    .X(_08371_));
 sky130_fd_sc_hd__mux2_1 _14782_ (.A0(\core.cpuregs[26][12] ),
    .A1(\core.cpuregs[27][12] ),
    .S(_08230_),
    .X(_08372_));
 sky130_fd_sc_hd__mux2_1 _14783_ (.A0(_08371_),
    .A1(_08372_),
    .S(_08226_),
    .X(_08373_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(\core.cpuregs[28][12] ),
    .A1(\core.cpuregs[29][12] ),
    .S(_08224_),
    .X(_08374_));
 sky130_fd_sc_hd__mux2_1 _14785_ (.A0(\core.cpuregs[30][12] ),
    .A1(\core.cpuregs[31][12] ),
    .S(_08234_),
    .X(_08375_));
 sky130_fd_sc_hd__mux2_1 _14786_ (.A0(_08374_),
    .A1(_08375_),
    .S(_08253_),
    .X(_08376_));
 sky130_fd_sc_hd__mux2_1 _14787_ (.A0(_08373_),
    .A1(_08376_),
    .S(_08238_),
    .X(_08377_));
 sky130_fd_sc_hd__mux2_1 _14788_ (.A0(_08370_),
    .A1(_08377_),
    .S(_08240_),
    .X(_08378_));
 sky130_fd_sc_hd__mux2_1 _14789_ (.A0(\core.cpuregs[0][12] ),
    .A1(\core.cpuregs[1][12] ),
    .S(_08224_),
    .X(_08379_));
 sky130_fd_sc_hd__mux2_4 _14790_ (.A0(\core.cpuregs[2][12] ),
    .A1(\core.cpuregs[3][12] ),
    .S(_06240_),
    .X(_08380_));
 sky130_fd_sc_hd__mux2_1 _14791_ (.A0(_08379_),
    .A1(_08380_),
    .S(_08226_),
    .X(_08381_));
 sky130_fd_sc_hd__mux2_1 _14792_ (.A0(\core.cpuregs[6][12] ),
    .A1(\core.cpuregs[7][12] ),
    .S(_08230_),
    .X(_08382_));
 sky130_fd_sc_hd__mux2_4 _14793_ (.A0(\core.cpuregs[4][12] ),
    .A1(\core.cpuregs[5][12] ),
    .S(_06256_),
    .X(_08383_));
 sky130_fd_sc_hd__mux2_1 _14794_ (.A0(_08382_),
    .A1(_08383_),
    .S(_08257_),
    .X(_08384_));
 sky130_fd_sc_hd__mux2_1 _14795_ (.A0(_08381_),
    .A1(_08384_),
    .S(_08249_),
    .X(_08385_));
 sky130_fd_sc_hd__mux2_1 _14796_ (.A0(\core.cpuregs[16][12] ),
    .A1(\core.cpuregs[17][12] ),
    .S(_08230_),
    .X(_08386_));
 sky130_fd_sc_hd__mux2_1 _14797_ (.A0(\core.cpuregs[18][12] ),
    .A1(\core.cpuregs[19][12] ),
    .S(_06256_),
    .X(_08387_));
 sky130_fd_sc_hd__mux2_1 _14798_ (.A0(_08386_),
    .A1(_08387_),
    .S(_08253_),
    .X(_08388_));
 sky130_fd_sc_hd__mux2_1 _14799_ (.A0(\core.cpuregs[22][12] ),
    .A1(\core.cpuregs[23][12] ),
    .S(_08234_),
    .X(_08389_));
 sky130_fd_sc_hd__mux2_4 _14800_ (.A0(\core.cpuregs[20][12] ),
    .A1(\core.cpuregs[21][12] ),
    .S(_06260_),
    .X(_08390_));
 sky130_fd_sc_hd__mux2_1 _14801_ (.A0(_08389_),
    .A1(_08390_),
    .S(_08257_),
    .X(_08391_));
 sky130_fd_sc_hd__mux2_4 _14802_ (.A0(_08388_),
    .A1(_08391_),
    .S(_08249_),
    .X(_08392_));
 sky130_fd_sc_hd__mux2_1 _14803_ (.A0(_08385_),
    .A1(_08392_),
    .S(_06268_),
    .X(_08393_));
 sky130_fd_sc_hd__mux2_1 _14804_ (.A0(_08378_),
    .A1(_08393_),
    .S(_06293_),
    .X(_08394_));
 sky130_fd_sc_hd__nand2_1 _14805_ (.A(_08394_),
    .B(_07722_),
    .Y(_08395_));
 sky130_fd_sc_hd__inv_2 _14806_ (.A(\core.reg_pc[12] ),
    .Y(_08396_));
 sky130_fd_sc_hd__or3_1 _14807_ (.A(_06302_),
    .B(_08396_),
    .C(_06305_),
    .X(_08397_));
 sky130_fd_sc_hd__a21o_1 _14808_ (.A1(_08395_),
    .A2(_08397_),
    .B1(_07894_),
    .X(_08398_));
 sky130_fd_sc_hd__a31o_1 _14809_ (.A1(_06099_),
    .A2(_06130_),
    .A3(_06138_),
    .B1(_06143_),
    .X(_08399_));
 sky130_fd_sc_hd__or2_1 _14810_ (.A(_06102_),
    .B(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_1 _14811_ (.A(_08399_),
    .B(_06102_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand3_1 _14812_ (.A(_08400_),
    .B(_06226_),
    .C(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__nand2_1 _14813_ (.A(_08270_),
    .B(_04792_),
    .Y(_08403_));
 sky130_fd_sc_hd__a21oi_2 _14814_ (.A1(_08403_),
    .A2(_08208_),
    .B1(_08272_),
    .Y(_08404_));
 sky130_fd_sc_hd__nand2_1 _14815_ (.A(_08117_),
    .B(_04901_),
    .Y(_08405_));
 sky130_fd_sc_hd__a21oi_1 _14816_ (.A1(_08206_),
    .A2(_08405_),
    .B1(_04589_),
    .Y(_08406_));
 sky130_fd_sc_hd__o31a_1 _14817_ (.A1(_04588_),
    .A2(_08404_),
    .A3(_08406_),
    .B1(_07651_),
    .X(_08407_));
 sky130_fd_sc_hd__nand3_1 _14818_ (.A(_08398_),
    .B(_08402_),
    .C(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand2_1 _14819_ (.A(_07728_),
    .B(_04796_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand2_1 _14820_ (.A(_08408_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__inv_2 _14821_ (.A(_08410_),
    .Y(_00255_));
 sky130_fd_sc_hd__mux2_1 _14822_ (.A0(\core.cpuregs[12][13] ),
    .A1(\core.cpuregs[13][13] ),
    .S(_08281_),
    .X(_08411_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(\core.cpuregs[14][13] ),
    .A1(\core.cpuregs[15][13] ),
    .S(_08283_),
    .X(_08412_));
 sky130_fd_sc_hd__mux2_1 _14824_ (.A0(_08411_),
    .A1(_08412_),
    .S(_08286_),
    .X(_08413_));
 sky130_fd_sc_hd__mux2_1 _14825_ (.A0(\core.cpuregs[8][13] ),
    .A1(\core.cpuregs[9][13] ),
    .S(_08288_),
    .X(_08414_));
 sky130_fd_sc_hd__mux2_1 _14826_ (.A0(\core.cpuregs[10][13] ),
    .A1(\core.cpuregs[11][13] ),
    .S(_08291_),
    .X(_08415_));
 sky130_fd_sc_hd__mux2_1 _14827_ (.A0(_08414_),
    .A1(_08415_),
    .S(_08294_),
    .X(_08416_));
 sky130_fd_sc_hd__clkbuf_2 _14828_ (.A(_06253_),
    .X(_08417_));
 sky130_fd_sc_hd__mux2_1 _14829_ (.A0(_08413_),
    .A1(_08416_),
    .S(_08417_),
    .X(_08418_));
 sky130_fd_sc_hd__mux2_1 _14830_ (.A0(\core.cpuregs[24][13] ),
    .A1(\core.cpuregs[25][13] ),
    .S(_08298_),
    .X(_08419_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(\core.cpuregs[26][13] ),
    .A1(\core.cpuregs[27][13] ),
    .S(_08300_),
    .X(_08420_));
 sky130_fd_sc_hd__mux2_1 _14832_ (.A0(_08419_),
    .A1(_08420_),
    .S(_08302_),
    .X(_08421_));
 sky130_fd_sc_hd__buf_4 _14833_ (.A(_08290_),
    .X(_08422_));
 sky130_fd_sc_hd__mux2_2 _14834_ (.A0(\core.cpuregs[28][13] ),
    .A1(\core.cpuregs[29][13] ),
    .S(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__clkbuf_4 _14835_ (.A(_08306_),
    .X(_08424_));
 sky130_fd_sc_hd__mux2_2 _14836_ (.A0(\core.cpuregs[30][13] ),
    .A1(\core.cpuregs[31][13] ),
    .S(_08424_),
    .X(_08425_));
 sky130_fd_sc_hd__mux2_1 _14837_ (.A0(_08423_),
    .A1(_08425_),
    .S(_08309_),
    .X(_08426_));
 sky130_fd_sc_hd__mux2_8 _14838_ (.A0(_08421_),
    .A1(_08426_),
    .S(_08311_),
    .X(_08427_));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(_08418_),
    .A1(_08427_),
    .S(_08313_),
    .X(_08428_));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(\core.cpuregs[0][13] ),
    .A1(\core.cpuregs[1][13] ),
    .S(_08315_),
    .X(_08429_));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(\core.cpuregs[2][13] ),
    .A1(\core.cpuregs[3][13] ),
    .S(_08317_),
    .X(_08430_));
 sky130_fd_sc_hd__mux2_1 _14842_ (.A0(_08429_),
    .A1(_08430_),
    .S(_08319_),
    .X(_08431_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(\core.cpuregs[6][13] ),
    .A1(\core.cpuregs[7][13] ),
    .S(_08321_),
    .X(_08432_));
 sky130_fd_sc_hd__mux2_1 _14844_ (.A0(\core.cpuregs[4][13] ),
    .A1(\core.cpuregs[5][13] ),
    .S(_08323_),
    .X(_08433_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(_08432_),
    .A1(_08433_),
    .S(_08325_),
    .X(_08434_));
 sky130_fd_sc_hd__mux2_2 _14846_ (.A0(_08431_),
    .A1(_08434_),
    .S(_08327_),
    .X(_08435_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\core.cpuregs[16][13] ),
    .A1(\core.cpuregs[17][13] ),
    .S(_08329_),
    .X(_08436_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(\core.cpuregs[18][13] ),
    .A1(\core.cpuregs[19][13] ),
    .S(_08323_),
    .X(_08437_));
 sky130_fd_sc_hd__clkbuf_4 _14849_ (.A(_08293_),
    .X(_08438_));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(_08436_),
    .A1(_08437_),
    .S(_08438_),
    .X(_08439_));
 sky130_fd_sc_hd__mux2_2 _14851_ (.A0(\core.cpuregs[22][13] ),
    .A1(\core.cpuregs[23][13] ),
    .S(_08334_),
    .X(_08440_));
 sky130_fd_sc_hd__mux2_1 _14852_ (.A0(\core.cpuregs[20][13] ),
    .A1(\core.cpuregs[21][13] ),
    .S(_08337_),
    .X(_08441_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(_08440_),
    .A1(_08441_),
    .S(_08339_),
    .X(_08442_));
 sky130_fd_sc_hd__mux2_1 _14854_ (.A0(_08439_),
    .A1(_08442_),
    .S(_08341_),
    .X(_08443_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(_08435_),
    .A1(_08443_),
    .S(_08343_),
    .X(_08444_));
 sky130_fd_sc_hd__mux2_1 _14856_ (.A0(_08428_),
    .A1(_08444_),
    .S(_08200_),
    .X(_08445_));
 sky130_fd_sc_hd__nand2_1 _14857_ (.A(_08445_),
    .B(_08202_),
    .Y(_08446_));
 sky130_fd_sc_hd__inv_2 _14858_ (.A(\core.reg_pc[13] ),
    .Y(_08447_));
 sky130_fd_sc_hd__or3_1 _14859_ (.A(_08347_),
    .B(_08447_),
    .C(_07852_),
    .X(_08448_));
 sky130_fd_sc_hd__nand2_1 _14860_ (.A(_08446_),
    .B(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__nand2_1 _14861_ (.A(_08449_),
    .B(_07783_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand2_1 _14862_ (.A(_08401_),
    .B(_06101_),
    .Y(_08451_));
 sky130_fd_sc_hd__a21oi_1 _14863_ (.A1(_08451_),
    .A2(_06105_),
    .B1(_04984_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21ai_1 _14864_ (.A1(_06105_),
    .A2(_08451_),
    .B1(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _14865_ (.A(_07790_),
    .B(_04796_),
    .Y(_08454_));
 sky130_fd_sc_hd__and3_1 _14866_ (.A(_08454_),
    .B(_08356_),
    .C(_08274_),
    .X(_08455_));
 sky130_fd_sc_hd__clkbuf_2 _14867_ (.A(_07786_),
    .X(_08456_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(_07901_),
    .B(_04904_),
    .Y(_08457_));
 sky130_fd_sc_hd__and3_1 _14869_ (.A(_08456_),
    .B(_08271_),
    .C(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__o21ai_1 _14870_ (.A1(_08455_),
    .A2(_08458_),
    .B1(_04634_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand3_2 _14871_ (.A(_08450_),
    .B(_08453_),
    .C(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_1 _14872_ (.A(_08460_),
    .B(_08215_),
    .Y(_08461_));
 sky130_fd_sc_hd__o21ai_1 _14873_ (.A1(_04799_),
    .A2(_08033_),
    .B1(_08461_),
    .Y(_00256_));
 sky130_fd_sc_hd__clkbuf_2 _14874_ (.A(_07651_),
    .X(_08462_));
 sky130_fd_sc_hd__mux2_1 _14875_ (.A0(\core.cpuregs[12][14] ),
    .A1(\core.cpuregs[13][14] ),
    .S(_08281_),
    .X(_08463_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(\core.cpuregs[14][14] ),
    .A1(\core.cpuregs[15][14] ),
    .S(_08283_),
    .X(_08464_));
 sky130_fd_sc_hd__mux2_1 _14877_ (.A0(_08463_),
    .A1(_08464_),
    .S(_08286_),
    .X(_08465_));
 sky130_fd_sc_hd__mux2_1 _14878_ (.A0(\core.cpuregs[8][14] ),
    .A1(\core.cpuregs[9][14] ),
    .S(_08288_),
    .X(_08466_));
 sky130_fd_sc_hd__mux2_1 _14879_ (.A0(\core.cpuregs[10][14] ),
    .A1(\core.cpuregs[11][14] ),
    .S(_08291_),
    .X(_08467_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(_08466_),
    .A1(_08467_),
    .S(_08294_),
    .X(_08468_));
 sky130_fd_sc_hd__mux2_1 _14881_ (.A0(_08465_),
    .A1(_08468_),
    .S(_08417_),
    .X(_08469_));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(\core.cpuregs[24][14] ),
    .A1(\core.cpuregs[25][14] ),
    .S(_08298_),
    .X(_08470_));
 sky130_fd_sc_hd__mux2_1 _14883_ (.A0(\core.cpuregs[26][14] ),
    .A1(\core.cpuregs[27][14] ),
    .S(_08300_),
    .X(_08471_));
 sky130_fd_sc_hd__mux2_1 _14884_ (.A0(_08470_),
    .A1(_08471_),
    .S(_08302_),
    .X(_08472_));
 sky130_fd_sc_hd__mux2_1 _14885_ (.A0(\core.cpuregs[28][14] ),
    .A1(\core.cpuregs[29][14] ),
    .S(_08422_),
    .X(_08473_));
 sky130_fd_sc_hd__mux2_1 _14886_ (.A0(\core.cpuregs[30][14] ),
    .A1(\core.cpuregs[31][14] ),
    .S(_08424_),
    .X(_08474_));
 sky130_fd_sc_hd__mux2_1 _14887_ (.A0(_08473_),
    .A1(_08474_),
    .S(_08332_),
    .X(_08475_));
 sky130_fd_sc_hd__mux2_1 _14888_ (.A0(_08472_),
    .A1(_08475_),
    .S(_08311_),
    .X(_08476_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(_08469_),
    .A1(_08476_),
    .S(_08313_),
    .X(_08477_));
 sky130_fd_sc_hd__mux2_1 _14890_ (.A0(\core.cpuregs[0][14] ),
    .A1(\core.cpuregs[1][14] ),
    .S(_08304_),
    .X(_08478_));
 sky130_fd_sc_hd__mux2_1 _14891_ (.A0(\core.cpuregs[2][14] ),
    .A1(\core.cpuregs[3][14] ),
    .S(_08307_),
    .X(_08479_));
 sky130_fd_sc_hd__mux2_1 _14892_ (.A0(_08478_),
    .A1(_08479_),
    .S(_08319_),
    .X(_08480_));
 sky130_fd_sc_hd__mux2_1 _14893_ (.A0(\core.cpuregs[6][14] ),
    .A1(\core.cpuregs[7][14] ),
    .S(_08321_),
    .X(_08481_));
 sky130_fd_sc_hd__buf_4 _14894_ (.A(_08336_),
    .X(_08482_));
 sky130_fd_sc_hd__mux2_1 _14895_ (.A0(\core.cpuregs[4][14] ),
    .A1(\core.cpuregs[5][14] ),
    .S(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__mux2_1 _14896_ (.A0(_08481_),
    .A1(_08483_),
    .S(_08325_),
    .X(_08484_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(_08480_),
    .A1(_08484_),
    .S(_08327_),
    .X(_08485_));
 sky130_fd_sc_hd__mux2_1 _14898_ (.A0(\core.cpuregs[16][14] ),
    .A1(\core.cpuregs[17][14] ),
    .S(_08329_),
    .X(_08486_));
 sky130_fd_sc_hd__mux2_1 _14899_ (.A0(\core.cpuregs[18][14] ),
    .A1(\core.cpuregs[19][14] ),
    .S(_08323_),
    .X(_08487_));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(_08486_),
    .A1(_08487_),
    .S(_08438_),
    .X(_08488_));
 sky130_fd_sc_hd__mux2_1 _14901_ (.A0(\core.cpuregs[22][14] ),
    .A1(\core.cpuregs[23][14] ),
    .S(_08334_),
    .X(_08489_));
 sky130_fd_sc_hd__mux2_1 _14902_ (.A0(\core.cpuregs[20][14] ),
    .A1(\core.cpuregs[21][14] ),
    .S(_08337_),
    .X(_08490_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(_08489_),
    .A1(_08490_),
    .S(_08339_),
    .X(_08491_));
 sky130_fd_sc_hd__mux2_1 _14904_ (.A0(_08488_),
    .A1(_08491_),
    .S(_08341_),
    .X(_08492_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(_08485_),
    .A1(_08492_),
    .S(_08343_),
    .X(_08493_));
 sky130_fd_sc_hd__mux2_1 _14906_ (.A0(_08477_),
    .A1(_08493_),
    .S(_08200_),
    .X(_08494_));
 sky130_fd_sc_hd__nand2_1 _14907_ (.A(_08494_),
    .B(_08202_),
    .Y(_08495_));
 sky130_fd_sc_hd__buf_2 _14908_ (.A(_06304_),
    .X(_08496_));
 sky130_fd_sc_hd__or3b_1 _14909_ (.A(_08347_),
    .B(_08496_),
    .C_N(_07355_),
    .X(_08497_));
 sky130_fd_sc_hd__nand2_1 _14910_ (.A(_08495_),
    .B(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__nand2_1 _14911_ (.A(_08498_),
    .B(_07783_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand2_1 _14912_ (.A(_08399_),
    .B(_06107_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_1 _14913_ (.A(_08500_),
    .B(_06144_),
    .Y(_08501_));
 sky130_fd_sc_hd__or2_1 _14914_ (.A(_06116_),
    .B(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__clkbuf_4 _14915_ (.A(_06225_),
    .X(_08503_));
 sky130_fd_sc_hd__nand2_1 _14916_ (.A(_08501_),
    .B(_06116_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand3_1 _14917_ (.A(_08502_),
    .B(_08503_),
    .C(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(_07657_),
    .B(_04799_),
    .Y(_08506_));
 sky130_fd_sc_hd__and3_1 _14919_ (.A(_08506_),
    .B(_08356_),
    .C(_08359_),
    .X(_08507_));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(_08358_),
    .B(_04909_),
    .Y(_08508_));
 sky130_fd_sc_hd__and3_1 _14921_ (.A(_08456_),
    .B(_08355_),
    .C(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__buf_1 _14922_ (.A(_04633_),
    .X(_08510_));
 sky130_fd_sc_hd__o21ai_1 _14923_ (.A1(_08507_),
    .A2(_08509_),
    .B1(_08510_),
    .Y(_08511_));
 sky130_fd_sc_hd__nand3_1 _14924_ (.A(_08499_),
    .B(_08505_),
    .C(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand2_1 _14925_ (.A(_08512_),
    .B(_08215_),
    .Y(_08513_));
 sky130_fd_sc_hd__o21ai_2 _14926_ (.A1(_04804_),
    .A2(_08462_),
    .B1(_08513_),
    .Y(_00257_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _14927_ (.A(_07682_),
    .X(_08514_));
 sky130_fd_sc_hd__buf_4 _14928_ (.A(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__mux2_1 _14929_ (.A0(\core.cpuregs[12][15] ),
    .A1(\core.cpuregs[13][15] ),
    .S(_08515_),
    .X(_08516_));
 sky130_fd_sc_hd__clkbuf_2 _14930_ (.A(_08514_),
    .X(_08517_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(\core.cpuregs[14][15] ),
    .A1(\core.cpuregs[15][15] ),
    .S(_08517_),
    .X(_08518_));
 sky130_fd_sc_hd__clkbuf_4 _14932_ (.A(_08285_),
    .X(_08519_));
 sky130_fd_sc_hd__mux2_1 _14933_ (.A0(_08516_),
    .A1(_08518_),
    .S(_08519_),
    .X(_08520_));
 sky130_fd_sc_hd__mux2_1 _14934_ (.A0(\core.cpuregs[8][15] ),
    .A1(\core.cpuregs[9][15] ),
    .S(_08517_),
    .X(_08521_));
 sky130_fd_sc_hd__clkbuf_2 _14935_ (.A(_08514_),
    .X(_08522_));
 sky130_fd_sc_hd__mux2_1 _14936_ (.A0(\core.cpuregs[10][15] ),
    .A1(\core.cpuregs[11][15] ),
    .S(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__clkbuf_2 _14937_ (.A(_08285_),
    .X(_08524_));
 sky130_fd_sc_hd__mux2_1 _14938_ (.A0(_08521_),
    .A1(_08523_),
    .S(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__mux2_1 _14939_ (.A0(_08520_),
    .A1(_08525_),
    .S(_08296_),
    .X(_08526_));
 sky130_fd_sc_hd__clkbuf_2 _14940_ (.A(_08514_),
    .X(_08527_));
 sky130_fd_sc_hd__mux2_1 _14941_ (.A0(\core.cpuregs[0][15] ),
    .A1(\core.cpuregs[1][15] ),
    .S(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__clkbuf_2 _14942_ (.A(_08280_),
    .X(_08529_));
 sky130_fd_sc_hd__mux2_1 _14943_ (.A0(\core.cpuregs[2][15] ),
    .A1(\core.cpuregs[3][15] ),
    .S(_08529_),
    .X(_08530_));
 sky130_fd_sc_hd__clkbuf_2 _14944_ (.A(_08285_),
    .X(_08531_));
 sky130_fd_sc_hd__mux2_1 _14945_ (.A0(_08528_),
    .A1(_08530_),
    .S(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__clkbuf_2 _14946_ (.A(_08514_),
    .X(_08533_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(\core.cpuregs[6][15] ),
    .A1(\core.cpuregs[7][15] ),
    .S(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__clkbuf_2 _14948_ (.A(_08280_),
    .X(_08535_));
 sky130_fd_sc_hd__mux2_2 _14949_ (.A0(\core.cpuregs[4][15] ),
    .A1(\core.cpuregs[5][15] ),
    .S(_08535_),
    .X(_08536_));
 sky130_fd_sc_hd__buf_4 _14950_ (.A(_07687_),
    .X(_08537_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(_08534_),
    .A1(_08536_),
    .S(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__clkbuf_2 _14952_ (.A(_07827_),
    .X(_08539_));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(_08532_),
    .A1(_08538_),
    .S(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__clkbuf_2 _14954_ (.A(_06291_),
    .X(_08541_));
 sky130_fd_sc_hd__mux2_1 _14955_ (.A0(_08526_),
    .A1(_08540_),
    .S(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__nand2_1 _14956_ (.A(_08542_),
    .B(_07848_),
    .Y(_08543_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(\core.cpuregs[24][15] ),
    .A1(\core.cpuregs[25][15] ),
    .S(_06240_),
    .X(_08544_));
 sky130_fd_sc_hd__mux2_1 _14958_ (.A0(\core.cpuregs[26][15] ),
    .A1(\core.cpuregs[27][15] ),
    .S(_06243_),
    .X(_08545_));
 sky130_fd_sc_hd__mux2_1 _14959_ (.A0(_08544_),
    .A1(_08545_),
    .S(_08253_),
    .X(_08546_));
 sky130_fd_sc_hd__mux2_4 _14960_ (.A0(\core.cpuregs[28][15] ),
    .A1(\core.cpuregs[29][15] ),
    .S(_06256_),
    .X(_08547_));
 sky130_fd_sc_hd__mux2_1 _14961_ (.A0(\core.cpuregs[30][15] ),
    .A1(\core.cpuregs[31][15] ),
    .S(_06250_),
    .X(_08548_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(_08547_),
    .A1(_08548_),
    .S(_06247_),
    .X(_08549_));
 sky130_fd_sc_hd__mux2_1 _14963_ (.A0(_08546_),
    .A1(_08549_),
    .S(_08249_),
    .X(_08550_));
 sky130_fd_sc_hd__mux2_2 _14964_ (.A0(\core.cpuregs[16][15] ),
    .A1(\core.cpuregs[17][15] ),
    .S(_06243_),
    .X(_08551_));
 sky130_fd_sc_hd__mux2_1 _14965_ (.A0(\core.cpuregs[18][15] ),
    .A1(\core.cpuregs[19][15] ),
    .S(_06273_),
    .X(_08552_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(_08551_),
    .A1(_08552_),
    .S(_06264_),
    .X(_08553_));
 sky130_fd_sc_hd__mux2_1 _14967_ (.A0(\core.cpuregs[22][15] ),
    .A1(\core.cpuregs[23][15] ),
    .S(_06250_),
    .X(_08554_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(\core.cpuregs[20][15] ),
    .A1(\core.cpuregs[21][15] ),
    .S(_06262_),
    .X(_08555_));
 sky130_fd_sc_hd__mux2_1 _14969_ (.A0(_08554_),
    .A1(_08555_),
    .S(_08257_),
    .X(_08556_));
 sky130_fd_sc_hd__mux2_1 _14970_ (.A0(_08553_),
    .A1(_08556_),
    .S(_06266_),
    .X(_08557_));
 sky130_fd_sc_hd__clkbuf_2 _14971_ (.A(_06291_),
    .X(_08558_));
 sky130_fd_sc_hd__mux2_1 _14972_ (.A0(_08550_),
    .A1(_08557_),
    .S(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__nand2_1 _14973_ (.A(_08559_),
    .B(_07720_),
    .Y(_08560_));
 sky130_fd_sc_hd__buf_4 _14974_ (.A(_06298_),
    .X(_08561_));
 sky130_fd_sc_hd__a21o_1 _14975_ (.A1(_08543_),
    .A2(_08560_),
    .B1(_08561_),
    .X(_08562_));
 sky130_fd_sc_hd__buf_1 _14976_ (.A(_06301_),
    .X(_08563_));
 sky130_fd_sc_hd__or3b_1 _14977_ (.A(_08563_),
    .B(_08065_),
    .C_N(_05275_),
    .X(_08564_));
 sky130_fd_sc_hd__a21o_1 _14978_ (.A1(_08562_),
    .A2(_08564_),
    .B1(_07894_),
    .X(_08565_));
 sky130_fd_sc_hd__nand2_1 _14979_ (.A(_08504_),
    .B(_06114_),
    .Y(_08566_));
 sky130_fd_sc_hd__or2_1 _14980_ (.A(_06111_),
    .B(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__nand2_1 _14981_ (.A(_08566_),
    .B(_06111_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand3_1 _14982_ (.A(_08567_),
    .B(_08503_),
    .C(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2_8 _14983_ (.A(_07657_),
    .B(_04804_),
    .Y(_08570_));
 sky130_fd_sc_hd__buf_1 _14984_ (.A(_07902_),
    .X(_08571_));
 sky130_fd_sc_hd__and3_1 _14985_ (.A(_08570_),
    .B(_08571_),
    .C(_08405_),
    .X(_08572_));
 sky130_fd_sc_hd__nand2_1 _14986_ (.A(_08358_),
    .B(_04911_),
    .Y(_08573_));
 sky130_fd_sc_hd__and3_1 _14987_ (.A(_08456_),
    .B(_08403_),
    .C(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__o21ai_1 _14988_ (.A1(_08572_),
    .A2(_08574_),
    .B1(_08510_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand3_1 _14989_ (.A(_08565_),
    .B(_08569_),
    .C(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_1 _14990_ (.A(_08576_),
    .B(_08215_),
    .Y(_08577_));
 sky130_fd_sc_hd__o21ai_1 _14991_ (.A1(_04806_),
    .A2(_08462_),
    .B1(_08577_),
    .Y(_00258_));
 sky130_fd_sc_hd__mux2_1 _14992_ (.A0(\core.cpuregs[12][16] ),
    .A1(\core.cpuregs[13][16] ),
    .S(_07919_),
    .X(_08578_));
 sky130_fd_sc_hd__mux2_1 _14993_ (.A0(\core.cpuregs[14][16] ),
    .A1(\core.cpuregs[15][16] ),
    .S(_07934_),
    .X(_08579_));
 sky130_fd_sc_hd__mux2_1 _14994_ (.A0(_08578_),
    .A1(_08579_),
    .S(_07984_),
    .X(_08580_));
 sky130_fd_sc_hd__mux2_1 _14995_ (.A0(\core.cpuregs[8][16] ),
    .A1(\core.cpuregs[9][16] ),
    .S(_07909_),
    .X(_08581_));
 sky130_fd_sc_hd__mux2_1 _14996_ (.A0(\core.cpuregs[10][16] ),
    .A1(\core.cpuregs[11][16] ),
    .S(_07922_),
    .X(_08582_));
 sky130_fd_sc_hd__mux2_1 _14997_ (.A0(_08581_),
    .A1(_08582_),
    .S(_07938_),
    .X(_08583_));
 sky130_fd_sc_hd__mux2_1 _14998_ (.A0(_08580_),
    .A1(_08583_),
    .S(_07673_),
    .X(_08584_));
 sky130_fd_sc_hd__mux2_1 _14999_ (.A0(\core.cpuregs[24][16] ),
    .A1(\core.cpuregs[25][16] ),
    .S(_08083_),
    .X(_08585_));
 sky130_fd_sc_hd__mux2_1 _15000_ (.A0(\core.cpuregs[26][16] ),
    .A1(\core.cpuregs[27][16] ),
    .S(_07991_),
    .X(_08586_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(_08585_),
    .A1(_08586_),
    .S(_07916_),
    .X(_08587_));
 sky130_fd_sc_hd__mux2_1 _15002_ (.A0(\core.cpuregs[28][16] ),
    .A1(\core.cpuregs[29][16] ),
    .S(_07914_),
    .X(_08588_));
 sky130_fd_sc_hd__mux2_1 _15003_ (.A0(\core.cpuregs[30][16] ),
    .A1(\core.cpuregs[31][16] ),
    .S(_07953_),
    .X(_08589_));
 sky130_fd_sc_hd__mux2_1 _15004_ (.A0(_08588_),
    .A1(_08589_),
    .S(_07951_),
    .X(_08590_));
 sky130_fd_sc_hd__mux2_1 _15005_ (.A0(_08587_),
    .A1(_08590_),
    .S(_07945_),
    .X(_08591_));
 sky130_fd_sc_hd__mux2_1 _15006_ (.A0(_08584_),
    .A1(_08591_),
    .S(_07998_),
    .X(_08592_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(\core.cpuregs[0][16] ),
    .A1(\core.cpuregs[1][16] ),
    .S(_07926_),
    .X(_08593_));
 sky130_fd_sc_hd__mux2_1 _15008_ (.A0(\core.cpuregs[2][16] ),
    .A1(\core.cpuregs[3][16] ),
    .S(_07928_),
    .X(_08594_));
 sky130_fd_sc_hd__mux2_1 _15009_ (.A0(_08593_),
    .A1(_08594_),
    .S(_07930_),
    .X(_08595_));
 sky130_fd_sc_hd__mux2_1 _15010_ (.A0(\core.cpuregs[6][16] ),
    .A1(\core.cpuregs[7][16] ),
    .S(_07936_),
    .X(_08596_));
 sky130_fd_sc_hd__mux2_1 _15011_ (.A0(\core.cpuregs[4][16] ),
    .A1(\core.cpuregs[5][16] ),
    .S(_07955_),
    .X(_08597_));
 sky130_fd_sc_hd__mux2_1 _15012_ (.A0(_08596_),
    .A1(_08597_),
    .S(_07957_),
    .X(_08598_));
 sky130_fd_sc_hd__mux2_1 _15013_ (.A0(_08595_),
    .A1(_08598_),
    .S(_08006_),
    .X(_08599_));
 sky130_fd_sc_hd__mux2_1 _15014_ (.A0(\core.cpuregs[16][16] ),
    .A1(\core.cpuregs[17][16] ),
    .S(_07940_),
    .X(_08600_));
 sky130_fd_sc_hd__mux2_1 _15015_ (.A0(\core.cpuregs[18][16] ),
    .A1(\core.cpuregs[19][16] ),
    .S(_08009_),
    .X(_08601_));
 sky130_fd_sc_hd__mux2_1 _15016_ (.A0(_08600_),
    .A1(_08601_),
    .S(_07712_),
    .X(_08602_));
 sky130_fd_sc_hd__mux2_1 _15017_ (.A0(\core.cpuregs[22][16] ),
    .A1(\core.cpuregs[23][16] ),
    .S(_07949_),
    .X(_08603_));
 sky130_fd_sc_hd__mux2_1 _15018_ (.A0(\core.cpuregs[20][16] ),
    .A1(\core.cpuregs[21][16] ),
    .S(_07684_),
    .X(_08604_));
 sky130_fd_sc_hd__mux2_1 _15019_ (.A0(_08603_),
    .A1(_08604_),
    .S(_07688_),
    .X(_08605_));
 sky130_fd_sc_hd__clkbuf_2 _15020_ (.A(_07827_),
    .X(_08606_));
 sky130_fd_sc_hd__mux2_1 _15021_ (.A0(_08602_),
    .A1(_08605_),
    .S(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__mux2_1 _15022_ (.A0(_08599_),
    .A1(_08607_),
    .S(_08313_),
    .X(_08608_));
 sky130_fd_sc_hd__mux2_1 _15023_ (.A0(_08592_),
    .A1(_08608_),
    .S(_08200_),
    .X(_08609_));
 sky130_fd_sc_hd__inv_2 _15024_ (.A(\core.reg_pc[16] ),
    .Y(_08610_));
 sky130_fd_sc_hd__or3_1 _15025_ (.A(_06301_),
    .B(_08610_),
    .C(_08065_),
    .X(_08611_));
 sky130_fd_sc_hd__a21boi_1 _15026_ (.A1(_08609_),
    .A2(_08202_),
    .B1_N(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_07656_),
    .B(_04806_),
    .Y(_08613_));
 sky130_fd_sc_hd__a21oi_1 _15028_ (.A1(_08613_),
    .A2(_08457_),
    .B1(_07786_),
    .Y(_08614_));
 sky130_fd_sc_hd__nand2_1 _15029_ (.A(_07802_),
    .B(_04917_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21oi_1 _15030_ (.A1(_08454_),
    .A2(_08615_),
    .B1(_08356_),
    .Y(_08616_));
 sky130_fd_sc_hd__or2_1 _15031_ (.A(_06178_),
    .B(_06148_),
    .X(_08617_));
 sky130_fd_sc_hd__nand2_1 _15032_ (.A(_06148_),
    .B(_06178_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_1 _15033_ (.A(_08617_),
    .B(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__o32a_1 _15034_ (.A1(_06230_),
    .A2(_08614_),
    .A3(_08616_),
    .B1(_04983_),
    .B2(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__o21ai_1 _15035_ (.A1(_08169_),
    .A2(_08612_),
    .B1(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand2_1 _15036_ (.A(_08621_),
    .B(_08215_),
    .Y(_08622_));
 sky130_fd_sc_hd__o21ai_1 _15037_ (.A1(_04901_),
    .A2(_08462_),
    .B1(_08622_),
    .Y(_00259_));
 sky130_fd_sc_hd__mux2_1 _15038_ (.A0(\core.cpuregs[12][17] ),
    .A1(\core.cpuregs[13][17] ),
    .S(_08281_),
    .X(_08623_));
 sky130_fd_sc_hd__mux2_1 _15039_ (.A0(\core.cpuregs[14][17] ),
    .A1(\core.cpuregs[15][17] ),
    .S(_08315_),
    .X(_08624_));
 sky130_fd_sc_hd__mux2_1 _15040_ (.A0(_08623_),
    .A1(_08624_),
    .S(_08286_),
    .X(_08625_));
 sky130_fd_sc_hd__mux2_1 _15041_ (.A0(\core.cpuregs[8][17] ),
    .A1(\core.cpuregs[9][17] ),
    .S(_08288_),
    .X(_08626_));
 sky130_fd_sc_hd__mux2_1 _15042_ (.A0(\core.cpuregs[10][17] ),
    .A1(\core.cpuregs[11][17] ),
    .S(_08291_),
    .X(_08627_));
 sky130_fd_sc_hd__mux2_1 _15043_ (.A0(_08626_),
    .A1(_08627_),
    .S(_08294_),
    .X(_08628_));
 sky130_fd_sc_hd__mux2_1 _15044_ (.A0(_08625_),
    .A1(_08628_),
    .S(_08417_),
    .X(_08629_));
 sky130_fd_sc_hd__mux2_1 _15045_ (.A0(\core.cpuregs[24][17] ),
    .A1(\core.cpuregs[25][17] ),
    .S(_08298_),
    .X(_08630_));
 sky130_fd_sc_hd__mux2_1 _15046_ (.A0(\core.cpuregs[26][17] ),
    .A1(\core.cpuregs[27][17] ),
    .S(_08300_),
    .X(_08631_));
 sky130_fd_sc_hd__mux2_1 _15047_ (.A0(_08630_),
    .A1(_08631_),
    .S(_08302_),
    .X(_08632_));
 sky130_fd_sc_hd__mux2_1 _15048_ (.A0(\core.cpuregs[28][17] ),
    .A1(\core.cpuregs[29][17] ),
    .S(_08422_),
    .X(_08633_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(\core.cpuregs[30][17] ),
    .A1(\core.cpuregs[31][17] ),
    .S(_08424_),
    .X(_08634_));
 sky130_fd_sc_hd__mux2_1 _15050_ (.A0(_08633_),
    .A1(_08634_),
    .S(_08332_),
    .X(_08635_));
 sky130_fd_sc_hd__mux2_1 _15051_ (.A0(_08632_),
    .A1(_08635_),
    .S(_08311_),
    .X(_08636_));
 sky130_fd_sc_hd__mux2_1 _15052_ (.A0(_08629_),
    .A1(_08636_),
    .S(_08313_),
    .X(_08637_));
 sky130_fd_sc_hd__mux2_1 _15053_ (.A0(\core.cpuregs[0][17] ),
    .A1(\core.cpuregs[1][17] ),
    .S(_08304_),
    .X(_08638_));
 sky130_fd_sc_hd__mux2_1 _15054_ (.A0(\core.cpuregs[2][17] ),
    .A1(\core.cpuregs[3][17] ),
    .S(_08307_),
    .X(_08639_));
 sky130_fd_sc_hd__mux2_1 _15055_ (.A0(_08638_),
    .A1(_08639_),
    .S(_08309_),
    .X(_08640_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(\core.cpuregs[6][17] ),
    .A1(\core.cpuregs[7][17] ),
    .S(_08317_),
    .X(_08641_));
 sky130_fd_sc_hd__mux2_1 _15057_ (.A0(\core.cpuregs[4][17] ),
    .A1(\core.cpuregs[5][17] ),
    .S(_08482_),
    .X(_08642_));
 sky130_fd_sc_hd__mux2_1 _15058_ (.A0(_08641_),
    .A1(_08642_),
    .S(_08325_),
    .X(_08643_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(_08640_),
    .A1(_08643_),
    .S(_08327_),
    .X(_08644_));
 sky130_fd_sc_hd__mux2_1 _15060_ (.A0(\core.cpuregs[16][17] ),
    .A1(\core.cpuregs[17][17] ),
    .S(_08329_),
    .X(_08645_));
 sky130_fd_sc_hd__mux2_1 _15061_ (.A0(\core.cpuregs[18][17] ),
    .A1(\core.cpuregs[19][17] ),
    .S(_08482_),
    .X(_08646_));
 sky130_fd_sc_hd__mux2_1 _15062_ (.A0(_08645_),
    .A1(_08646_),
    .S(_08438_),
    .X(_08647_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(\core.cpuregs[22][17] ),
    .A1(\core.cpuregs[23][17] ),
    .S(_08334_),
    .X(_08648_));
 sky130_fd_sc_hd__buf_4 _15064_ (.A(_08336_),
    .X(_08649_));
 sky130_fd_sc_hd__mux2_1 _15065_ (.A0(\core.cpuregs[20][17] ),
    .A1(\core.cpuregs[21][17] ),
    .S(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__mux2_2 _15066_ (.A0(_08648_),
    .A1(_08650_),
    .S(_08339_),
    .X(_08651_));
 sky130_fd_sc_hd__clkbuf_2 _15067_ (.A(_08237_),
    .X(_08652_));
 sky130_fd_sc_hd__mux2_1 _15068_ (.A0(_08647_),
    .A1(_08651_),
    .S(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__mux2_1 _15069_ (.A0(_08644_),
    .A1(_08653_),
    .S(_08343_),
    .X(_08654_));
 sky130_fd_sc_hd__mux2_1 _15070_ (.A0(_08637_),
    .A1(_08654_),
    .S(_08200_),
    .X(_08655_));
 sky130_fd_sc_hd__nand2_1 _15071_ (.A(_08655_),
    .B(_08202_),
    .Y(_08656_));
 sky130_fd_sc_hd__inv_2 _15072_ (.A(\core.reg_pc[17] ),
    .Y(_08657_));
 sky130_fd_sc_hd__or3_1 _15073_ (.A(_08347_),
    .B(_08657_),
    .C(_06305_),
    .X(_08658_));
 sky130_fd_sc_hd__nand2_1 _15074_ (.A(_08656_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2_2 _15075_ (.A(_08659_),
    .B(_07783_),
    .Y(_08660_));
 sky130_fd_sc_hd__nand2_1 _15076_ (.A(_08618_),
    .B(_06177_),
    .Y(_08661_));
 sky130_fd_sc_hd__a21oi_1 _15077_ (.A1(_08661_),
    .A2(_06175_),
    .B1(_04984_),
    .Y(_08662_));
 sky130_fd_sc_hd__o21ai_2 _15078_ (.A1(_06175_),
    .A2(_08661_),
    .B1(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand2_1 _15079_ (.A(_07657_),
    .B(_04901_),
    .Y(_08664_));
 sky130_fd_sc_hd__and3_1 _15080_ (.A(_08664_),
    .B(_08571_),
    .C(_08508_),
    .X(_08665_));
 sky130_fd_sc_hd__nand2_2 _15081_ (.A(_08358_),
    .B(_04916_),
    .Y(_08666_));
 sky130_fd_sc_hd__and3_1 _15082_ (.A(_08456_),
    .B(_08506_),
    .C(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__o21ai_2 _15083_ (.A1(_08665_),
    .A2(_08667_),
    .B1(_08510_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand3_1 _15084_ (.A(_08660_),
    .B(_08663_),
    .C(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15085_ (.A(_07724_),
    .X(_08670_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(_08669_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__o21ai_2 _15087_ (.A1(_04904_),
    .A2(_08462_),
    .B1(_08671_),
    .Y(_00260_));
 sky130_fd_sc_hd__mux2_1 _15088_ (.A0(\core.cpuregs[12][18] ),
    .A1(\core.cpuregs[13][18] ),
    .S(_08281_),
    .X(_08672_));
 sky130_fd_sc_hd__mux2_1 _15089_ (.A0(\core.cpuregs[14][18] ),
    .A1(\core.cpuregs[15][18] ),
    .S(_08315_),
    .X(_08673_));
 sky130_fd_sc_hd__mux2_1 _15090_ (.A0(_08672_),
    .A1(_08673_),
    .S(_08286_),
    .X(_08674_));
 sky130_fd_sc_hd__mux2_1 _15091_ (.A0(\core.cpuregs[8][18] ),
    .A1(\core.cpuregs[9][18] ),
    .S(_08288_),
    .X(_08675_));
 sky130_fd_sc_hd__mux2_1 _15092_ (.A0(\core.cpuregs[10][18] ),
    .A1(\core.cpuregs[11][18] ),
    .S(_08291_),
    .X(_08676_));
 sky130_fd_sc_hd__mux2_1 _15093_ (.A0(_08675_),
    .A1(_08676_),
    .S(_08319_),
    .X(_08677_));
 sky130_fd_sc_hd__mux2_1 _15094_ (.A0(_08674_),
    .A1(_08677_),
    .S(_08417_),
    .X(_08678_));
 sky130_fd_sc_hd__mux2_1 _15095_ (.A0(\core.cpuregs[24][18] ),
    .A1(\core.cpuregs[25][18] ),
    .S(_08283_),
    .X(_08679_));
 sky130_fd_sc_hd__mux2_1 _15096_ (.A0(\core.cpuregs[26][18] ),
    .A1(\core.cpuregs[27][18] ),
    .S(_08300_),
    .X(_08680_));
 sky130_fd_sc_hd__mux2_1 _15097_ (.A0(_08679_),
    .A1(_08680_),
    .S(_08302_),
    .X(_08681_));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(\core.cpuregs[28][18] ),
    .A1(\core.cpuregs[29][18] ),
    .S(_08422_),
    .X(_08682_));
 sky130_fd_sc_hd__mux2_2 _15099_ (.A0(\core.cpuregs[30][18] ),
    .A1(\core.cpuregs[31][18] ),
    .S(_08424_),
    .X(_08683_));
 sky130_fd_sc_hd__mux2_1 _15100_ (.A0(_08682_),
    .A1(_08683_),
    .S(_08332_),
    .X(_08684_));
 sky130_fd_sc_hd__mux2_8 _15101_ (.A0(_08681_),
    .A1(_08684_),
    .S(_08311_),
    .X(_08685_));
 sky130_fd_sc_hd__mux2_1 _15102_ (.A0(_08678_),
    .A1(_08685_),
    .S(_08313_),
    .X(_08686_));
 sky130_fd_sc_hd__mux2_1 _15103_ (.A0(\core.cpuregs[0][18] ),
    .A1(\core.cpuregs[1][18] ),
    .S(_08304_),
    .X(_08687_));
 sky130_fd_sc_hd__mux2_2 _15104_ (.A0(\core.cpuregs[2][18] ),
    .A1(\core.cpuregs[3][18] ),
    .S(_08307_),
    .X(_08688_));
 sky130_fd_sc_hd__mux2_1 _15105_ (.A0(_08687_),
    .A1(_08688_),
    .S(_08309_),
    .X(_08689_));
 sky130_fd_sc_hd__mux2_1 _15106_ (.A0(\core.cpuregs[6][18] ),
    .A1(\core.cpuregs[7][18] ),
    .S(_08317_),
    .X(_08690_));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(\core.cpuregs[4][18] ),
    .A1(\core.cpuregs[5][18] ),
    .S(_08482_),
    .X(_08691_));
 sky130_fd_sc_hd__mux2_1 _15108_ (.A0(_08690_),
    .A1(_08691_),
    .S(_08325_),
    .X(_08692_));
 sky130_fd_sc_hd__mux2_1 _15109_ (.A0(_08689_),
    .A1(_08692_),
    .S(_08341_),
    .X(_08693_));
 sky130_fd_sc_hd__mux2_1 _15110_ (.A0(\core.cpuregs[16][18] ),
    .A1(\core.cpuregs[17][18] ),
    .S(_08321_),
    .X(_08694_));
 sky130_fd_sc_hd__mux2_1 _15111_ (.A0(\core.cpuregs[18][18] ),
    .A1(\core.cpuregs[19][18] ),
    .S(_08482_),
    .X(_08695_));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(_08694_),
    .A1(_08695_),
    .S(_08438_),
    .X(_08696_));
 sky130_fd_sc_hd__mux2_1 _15113_ (.A0(\core.cpuregs[22][18] ),
    .A1(\core.cpuregs[23][18] ),
    .S(_08334_),
    .X(_08697_));
 sky130_fd_sc_hd__mux2_1 _15114_ (.A0(\core.cpuregs[20][18] ),
    .A1(\core.cpuregs[21][18] ),
    .S(_08649_),
    .X(_08698_));
 sky130_fd_sc_hd__mux2_1 _15115_ (.A0(_08697_),
    .A1(_08698_),
    .S(_08339_),
    .X(_08699_));
 sky130_fd_sc_hd__mux2_1 _15116_ (.A0(_08696_),
    .A1(_08699_),
    .S(_08652_),
    .X(_08700_));
 sky130_fd_sc_hd__mux2_8 _15117_ (.A0(_08693_),
    .A1(_08700_),
    .S(_08240_),
    .X(_08701_));
 sky130_fd_sc_hd__mux2_1 _15118_ (.A0(_08686_),
    .A1(_08701_),
    .S(_06293_),
    .X(_08702_));
 sky130_fd_sc_hd__nand2_1 _15119_ (.A(_08702_),
    .B(_07722_),
    .Y(_08703_));
 sky130_fd_sc_hd__or3b_1 _15120_ (.A(_08347_),
    .B(_08496_),
    .C_N(_05339_),
    .X(_08704_));
 sky130_fd_sc_hd__nand2_1 _15121_ (.A(_08703_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__nand2_2 _15122_ (.A(_08705_),
    .B(_07783_),
    .Y(_08706_));
 sky130_fd_sc_hd__a21o_2 _15123_ (.A1(_06140_),
    .A2(_06147_),
    .B1(_06179_),
    .X(_08707_));
 sky130_fd_sc_hd__nand2_2 _15124_ (.A(_08707_),
    .B(_06184_),
    .Y(_08708_));
 sky130_fd_sc_hd__or2_1 _15125_ (.A(_06167_),
    .B(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__nand2_1 _15126_ (.A(_08708_),
    .B(_06167_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand3_1 _15127_ (.A(_08709_),
    .B(_08503_),
    .C(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_1 _15128_ (.A(_08270_),
    .B(_04904_),
    .Y(_08712_));
 sky130_fd_sc_hd__and3_1 _15129_ (.A(_08712_),
    .B(_08571_),
    .C(_08573_),
    .X(_08713_));
 sky130_fd_sc_hd__nand2_1 _15130_ (.A(_08358_),
    .B(_04924_),
    .Y(_08714_));
 sky130_fd_sc_hd__and3_1 _15131_ (.A(_08456_),
    .B(_08570_),
    .C(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__o21ai_1 _15132_ (.A1(_08713_),
    .A2(_08715_),
    .B1(_08510_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand3_2 _15133_ (.A(_08706_),
    .B(_08711_),
    .C(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nand2_1 _15134_ (.A(_08717_),
    .B(_08670_),
    .Y(_08718_));
 sky130_fd_sc_hd__o21ai_1 _15135_ (.A1(_04909_),
    .A2(_08462_),
    .B1(_08718_),
    .Y(_00261_));
 sky130_fd_sc_hd__mux2_1 _15136_ (.A0(\core.cpuregs[12][19] ),
    .A1(\core.cpuregs[13][19] ),
    .S(_07692_),
    .X(_08719_));
 sky130_fd_sc_hd__clkbuf_4 _15137_ (.A(_07691_),
    .X(_08720_));
 sky130_fd_sc_hd__mux2_1 _15138_ (.A0(\core.cpuregs[14][19] ),
    .A1(\core.cpuregs[15][19] ),
    .S(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__clkbuf_4 _15139_ (.A(_08285_),
    .X(_08722_));
 sky130_fd_sc_hd__mux2_1 _15140_ (.A0(_08719_),
    .A1(_08721_),
    .S(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__mux2_1 _15141_ (.A0(\core.cpuregs[8][19] ),
    .A1(\core.cpuregs[9][19] ),
    .S(_08720_),
    .X(_08724_));
 sky130_fd_sc_hd__clkbuf_4 _15142_ (.A(_07691_),
    .X(_08725_));
 sky130_fd_sc_hd__mux2_1 _15143_ (.A0(\core.cpuregs[10][19] ),
    .A1(\core.cpuregs[11][19] ),
    .S(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__mux2_1 _15144_ (.A0(_08724_),
    .A1(_08726_),
    .S(_08722_),
    .X(_08727_));
 sky130_fd_sc_hd__mux2_1 _15145_ (.A0(_08723_),
    .A1(_08727_),
    .S(_07696_),
    .X(_08728_));
 sky130_fd_sc_hd__mux2_1 _15146_ (.A0(\core.cpuregs[0][19] ),
    .A1(\core.cpuregs[1][19] ),
    .S(_08720_),
    .X(_08729_));
 sky130_fd_sc_hd__mux2_1 _15147_ (.A0(\core.cpuregs[2][19] ),
    .A1(\core.cpuregs[3][19] ),
    .S(_08725_),
    .X(_08730_));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(_08729_),
    .A1(_08730_),
    .S(_08722_),
    .X(_08731_));
 sky130_fd_sc_hd__mux2_1 _15149_ (.A0(\core.cpuregs[6][19] ),
    .A1(\core.cpuregs[7][19] ),
    .S(_08725_),
    .X(_08732_));
 sky130_fd_sc_hd__clkbuf_4 _15150_ (.A(_07691_),
    .X(_08733_));
 sky130_fd_sc_hd__mux2_1 _15151_ (.A0(\core.cpuregs[4][19] ),
    .A1(\core.cpuregs[5][19] ),
    .S(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__mux2_1 _15152_ (.A0(_08732_),
    .A1(_08734_),
    .S(_07694_),
    .X(_08735_));
 sky130_fd_sc_hd__mux2_1 _15153_ (.A0(_08731_),
    .A1(_08735_),
    .S(_08606_),
    .X(_08736_));
 sky130_fd_sc_hd__clkbuf_4 _15154_ (.A(_06291_),
    .X(_08737_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(_08728_),
    .A1(_08736_),
    .S(_08737_),
    .X(_08738_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15156_ (.A(_07757_),
    .X(_08739_));
 sky130_fd_sc_hd__nand2_1 _15157_ (.A(_08738_),
    .B(_08739_),
    .Y(_08740_));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(\core.cpuregs[24][19] ),
    .A1(\core.cpuregs[25][19] ),
    .S(_08515_),
    .X(_08741_));
 sky130_fd_sc_hd__mux2_1 _15159_ (.A0(\core.cpuregs[26][19] ),
    .A1(\core.cpuregs[27][19] ),
    .S(_08527_),
    .X(_08742_));
 sky130_fd_sc_hd__mux2_1 _15160_ (.A0(_08741_),
    .A1(_08742_),
    .S(_08524_),
    .X(_08743_));
 sky130_fd_sc_hd__mux2_1 _15161_ (.A0(\core.cpuregs[28][19] ),
    .A1(\core.cpuregs[29][19] ),
    .S(_08527_),
    .X(_08744_));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(\core.cpuregs[30][19] ),
    .A1(\core.cpuregs[31][19] ),
    .S(_08533_),
    .X(_08745_));
 sky130_fd_sc_hd__mux2_1 _15163_ (.A0(_08744_),
    .A1(_08745_),
    .S(_08524_),
    .X(_08746_));
 sky130_fd_sc_hd__mux2_1 _15164_ (.A0(_08743_),
    .A1(_08746_),
    .S(_08539_),
    .X(_08747_));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(\core.cpuregs[16][19] ),
    .A1(\core.cpuregs[17][19] ),
    .S(_08522_),
    .X(_08748_));
 sky130_fd_sc_hd__mux2_1 _15166_ (.A0(\core.cpuregs[18][19] ),
    .A1(\core.cpuregs[19][19] ),
    .S(_08529_),
    .X(_08749_));
 sky130_fd_sc_hd__mux2_1 _15167_ (.A0(_08748_),
    .A1(_08749_),
    .S(_08531_),
    .X(_08750_));
 sky130_fd_sc_hd__mux2_1 _15168_ (.A0(\core.cpuregs[22][19] ),
    .A1(\core.cpuregs[23][19] ),
    .S(_08529_),
    .X(_08751_));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(\core.cpuregs[20][19] ),
    .A1(\core.cpuregs[21][19] ),
    .S(_08535_),
    .X(_08752_));
 sky130_fd_sc_hd__mux2_1 _15170_ (.A0(_08751_),
    .A1(_08752_),
    .S(_08537_),
    .X(_08753_));
 sky130_fd_sc_hd__mux2_1 _15171_ (.A0(_08750_),
    .A1(_08753_),
    .S(_08539_),
    .X(_08754_));
 sky130_fd_sc_hd__mux2_1 _15172_ (.A0(_08747_),
    .A1(_08754_),
    .S(_08541_),
    .X(_08755_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15173_ (.A(_07719_),
    .X(_08756_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(_08755_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__a21o_1 _15175_ (.A1(_08740_),
    .A2(_08757_),
    .B1(_07760_),
    .X(_08758_));
 sky130_fd_sc_hd__inv_2 _15176_ (.A(\core.reg_pc[19] ),
    .Y(_08759_));
 sky130_fd_sc_hd__or3_2 _15177_ (.A(_06302_),
    .B(_08759_),
    .C(_08496_),
    .X(_08760_));
 sky130_fd_sc_hd__nand2_8 _15178_ (.A(_08758_),
    .B(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand2_1 _15179_ (.A(_07656_),
    .B(_04909_),
    .Y(_08762_));
 sky130_fd_sc_hd__and3_1 _15180_ (.A(_08762_),
    .B(_04626_),
    .C(_08615_),
    .X(_08763_));
 sky130_fd_sc_hd__nand2_1 _15181_ (.A(_07901_),
    .B(_04922_),
    .Y(_08764_));
 sky130_fd_sc_hd__and3_1 _15182_ (.A(_07786_),
    .B(_08613_),
    .C(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__o21a_1 _15183_ (.A1(_08763_),
    .A2(_08765_),
    .B1(_05199_),
    .X(_08766_));
 sky130_fd_sc_hd__a21oi_4 _15184_ (.A1(_08761_),
    .A2(_06309_),
    .B1(_08766_),
    .Y(_08767_));
 sky130_fd_sc_hd__nand2_1 _15185_ (.A(_08710_),
    .B(_06166_),
    .Y(_08768_));
 sky130_fd_sc_hd__a21oi_2 _15186_ (.A1(_08768_),
    .A2(_06171_),
    .B1(_04984_),
    .Y(_08769_));
 sky130_fd_sc_hd__o21ai_4 _15187_ (.A1(_06171_),
    .A2(_08768_),
    .B1(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__nand2_8 _15188_ (.A(_08767_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_1 _15189_ (.A(_08771_),
    .B(_08670_),
    .Y(_08772_));
 sky130_fd_sc_hd__o21ai_1 _15190_ (.A1(_04911_),
    .A2(_08462_),
    .B1(_08772_),
    .Y(_00262_));
 sky130_fd_sc_hd__clkbuf_2 _15191_ (.A(_07651_),
    .X(_08773_));
 sky130_fd_sc_hd__mux2_1 _15192_ (.A0(\core.cpuregs[12][20] ),
    .A1(\core.cpuregs[13][20] ),
    .S(_08281_),
    .X(_08774_));
 sky130_fd_sc_hd__mux2_1 _15193_ (.A0(\core.cpuregs[14][20] ),
    .A1(\core.cpuregs[15][20] ),
    .S(_08315_),
    .X(_08775_));
 sky130_fd_sc_hd__mux2_1 _15194_ (.A0(_08774_),
    .A1(_08775_),
    .S(_08286_),
    .X(_08776_));
 sky130_fd_sc_hd__mux2_1 _15195_ (.A0(\core.cpuregs[8][20] ),
    .A1(\core.cpuregs[9][20] ),
    .S(_08298_),
    .X(_08777_));
 sky130_fd_sc_hd__mux2_1 _15196_ (.A0(\core.cpuregs[10][20] ),
    .A1(\core.cpuregs[11][20] ),
    .S(_08291_),
    .X(_08778_));
 sky130_fd_sc_hd__mux2_1 _15197_ (.A0(_08777_),
    .A1(_08778_),
    .S(_08319_),
    .X(_08779_));
 sky130_fd_sc_hd__mux2_1 _15198_ (.A0(_08776_),
    .A1(_08779_),
    .S(_08417_),
    .X(_08780_));
 sky130_fd_sc_hd__mux2_1 _15199_ (.A0(\core.cpuregs[24][20] ),
    .A1(\core.cpuregs[25][20] ),
    .S(_08283_),
    .X(_08781_));
 sky130_fd_sc_hd__mux2_2 _15200_ (.A0(\core.cpuregs[26][20] ),
    .A1(\core.cpuregs[27][20] ),
    .S(_08329_),
    .X(_08782_));
 sky130_fd_sc_hd__mux2_1 _15201_ (.A0(_08781_),
    .A1(_08782_),
    .S(_08294_),
    .X(_08783_));
 sky130_fd_sc_hd__mux2_1 _15202_ (.A0(\core.cpuregs[28][20] ),
    .A1(\core.cpuregs[29][20] ),
    .S(_08422_),
    .X(_08784_));
 sky130_fd_sc_hd__mux2_1 _15203_ (.A0(\core.cpuregs[30][20] ),
    .A1(\core.cpuregs[31][20] ),
    .S(_08424_),
    .X(_08785_));
 sky130_fd_sc_hd__mux2_1 _15204_ (.A0(_08784_),
    .A1(_08785_),
    .S(_08332_),
    .X(_08786_));
 sky130_fd_sc_hd__mux2_1 _15205_ (.A0(_08783_),
    .A1(_08786_),
    .S(_08327_),
    .X(_08787_));
 sky130_fd_sc_hd__mux2_2 _15206_ (.A0(_08780_),
    .A1(_08787_),
    .S(_08343_),
    .X(_08788_));
 sky130_fd_sc_hd__mux2_1 _15207_ (.A0(\core.cpuregs[0][20] ),
    .A1(\core.cpuregs[1][20] ),
    .S(_08304_),
    .X(_08789_));
 sky130_fd_sc_hd__mux2_1 _15208_ (.A0(\core.cpuregs[2][20] ),
    .A1(\core.cpuregs[3][20] ),
    .S(_08307_),
    .X(_08790_));
 sky130_fd_sc_hd__mux2_1 _15209_ (.A0(_08789_),
    .A1(_08790_),
    .S(_08309_),
    .X(_08791_));
 sky130_fd_sc_hd__mux2_1 _15210_ (.A0(\core.cpuregs[6][20] ),
    .A1(\core.cpuregs[7][20] ),
    .S(_08317_),
    .X(_08792_));
 sky130_fd_sc_hd__mux2_2 _15211_ (.A0(\core.cpuregs[4][20] ),
    .A1(\core.cpuregs[5][20] ),
    .S(_08337_),
    .X(_08793_));
 sky130_fd_sc_hd__mux2_1 _15212_ (.A0(_08792_),
    .A1(_08793_),
    .S(_08325_),
    .X(_08794_));
 sky130_fd_sc_hd__mux2_1 _15213_ (.A0(_08791_),
    .A1(_08794_),
    .S(_08341_),
    .X(_08795_));
 sky130_fd_sc_hd__mux2_1 _15214_ (.A0(\core.cpuregs[16][20] ),
    .A1(\core.cpuregs[17][20] ),
    .S(_08321_),
    .X(_08796_));
 sky130_fd_sc_hd__mux2_1 _15215_ (.A0(\core.cpuregs[18][20] ),
    .A1(\core.cpuregs[19][20] ),
    .S(_08482_),
    .X(_08797_));
 sky130_fd_sc_hd__mux2_1 _15216_ (.A0(_08796_),
    .A1(_08797_),
    .S(_08438_),
    .X(_08798_));
 sky130_fd_sc_hd__mux2_1 _15217_ (.A0(\core.cpuregs[22][20] ),
    .A1(\core.cpuregs[23][20] ),
    .S(_08334_),
    .X(_08799_));
 sky130_fd_sc_hd__mux2_2 _15218_ (.A0(\core.cpuregs[20][20] ),
    .A1(\core.cpuregs[21][20] ),
    .S(_08649_),
    .X(_08800_));
 sky130_fd_sc_hd__mux2_1 _15219_ (.A0(_08799_),
    .A1(_08800_),
    .S(_08247_),
    .X(_08801_));
 sky130_fd_sc_hd__mux2_2 _15220_ (.A0(_08798_),
    .A1(_08801_),
    .S(_08652_),
    .X(_08802_));
 sky130_fd_sc_hd__mux2_1 _15221_ (.A0(_08795_),
    .A1(_08802_),
    .S(_08240_),
    .X(_08803_));
 sky130_fd_sc_hd__mux2_1 _15222_ (.A0(_08788_),
    .A1(_08803_),
    .S(_06293_),
    .X(_08804_));
 sky130_fd_sc_hd__nand2_1 _15223_ (.A(_08804_),
    .B(_07722_),
    .Y(_08805_));
 sky130_fd_sc_hd__inv_2 _15224_ (.A(\core.reg_pc[20] ),
    .Y(_08806_));
 sky130_fd_sc_hd__or3_1 _15225_ (.A(_08347_),
    .B(_08806_),
    .C(_06305_),
    .X(_08807_));
 sky130_fd_sc_hd__nand2_1 _15226_ (.A(_08805_),
    .B(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(_08808_),
    .B(_06309_),
    .Y(_08809_));
 sky130_fd_sc_hd__nand2_1 _15228_ (.A(_06148_),
    .B(_06180_),
    .Y(_08810_));
 sky130_fd_sc_hd__inv_2 _15229_ (.A(_06185_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_08810_),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__or2_1 _15231_ (.A(_06163_),
    .B(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__nand2_1 _15232_ (.A(_08812_),
    .B(_06163_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand3_1 _15233_ (.A(_08813_),
    .B(_08503_),
    .C(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_2 _15234_ (.A(_08270_),
    .B(_04911_),
    .Y(_08816_));
 sky130_fd_sc_hd__and3_1 _15235_ (.A(_08816_),
    .B(_08571_),
    .C(_08666_),
    .X(_08817_));
 sky130_fd_sc_hd__nand2_1 _15236_ (.A(_06235_),
    .B(_04939_),
    .Y(_08818_));
 sky130_fd_sc_hd__and3_1 _15237_ (.A(_08456_),
    .B(_08664_),
    .C(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__o21ai_1 _15238_ (.A1(_08817_),
    .A2(_08819_),
    .B1(_08510_),
    .Y(_08820_));
 sky130_fd_sc_hd__nand3_1 _15239_ (.A(_08809_),
    .B(_08815_),
    .C(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand2_1 _15240_ (.A(_08821_),
    .B(_08670_),
    .Y(_08822_));
 sky130_fd_sc_hd__o21ai_1 _15241_ (.A1(_04917_),
    .A2(_08773_),
    .B1(_08822_),
    .Y(_00263_));
 sky130_fd_sc_hd__mux2_1 _15242_ (.A0(\core.cpuregs[12][21] ),
    .A1(\core.cpuregs[13][21] ),
    .S(_08515_),
    .X(_08823_));
 sky130_fd_sc_hd__mux2_1 _15243_ (.A0(\core.cpuregs[14][21] ),
    .A1(\core.cpuregs[15][21] ),
    .S(_08517_),
    .X(_08824_));
 sky130_fd_sc_hd__mux2_1 _15244_ (.A0(_08823_),
    .A1(_08824_),
    .S(_08519_),
    .X(_08825_));
 sky130_fd_sc_hd__mux2_1 _15245_ (.A0(\core.cpuregs[8][21] ),
    .A1(\core.cpuregs[9][21] ),
    .S(_08517_),
    .X(_08826_));
 sky130_fd_sc_hd__mux2_1 _15246_ (.A0(\core.cpuregs[10][21] ),
    .A1(\core.cpuregs[11][21] ),
    .S(_08522_),
    .X(_08827_));
 sky130_fd_sc_hd__mux2_1 _15247_ (.A0(_08826_),
    .A1(_08827_),
    .S(_08524_),
    .X(_08828_));
 sky130_fd_sc_hd__mux2_1 _15248_ (.A0(_08825_),
    .A1(_08828_),
    .S(_08296_),
    .X(_08829_));
 sky130_fd_sc_hd__mux2_1 _15249_ (.A0(\core.cpuregs[0][21] ),
    .A1(\core.cpuregs[1][21] ),
    .S(_08522_),
    .X(_08830_));
 sky130_fd_sc_hd__mux2_1 _15250_ (.A0(\core.cpuregs[2][21] ),
    .A1(\core.cpuregs[3][21] ),
    .S(_08529_),
    .X(_08831_));
 sky130_fd_sc_hd__mux2_1 _15251_ (.A0(_08830_),
    .A1(_08831_),
    .S(_08531_),
    .X(_08832_));
 sky130_fd_sc_hd__mux2_1 _15252_ (.A0(\core.cpuregs[6][21] ),
    .A1(\core.cpuregs[7][21] ),
    .S(_08533_),
    .X(_08833_));
 sky130_fd_sc_hd__mux2_4 _15253_ (.A0(\core.cpuregs[4][21] ),
    .A1(\core.cpuregs[5][21] ),
    .S(_08535_),
    .X(_08834_));
 sky130_fd_sc_hd__mux2_1 _15254_ (.A0(_08833_),
    .A1(_08834_),
    .S(_08537_),
    .X(_08835_));
 sky130_fd_sc_hd__mux2_1 _15255_ (.A0(_08832_),
    .A1(_08835_),
    .S(_08539_),
    .X(_08836_));
 sky130_fd_sc_hd__mux2_1 _15256_ (.A0(_08829_),
    .A1(_08836_),
    .S(_08541_),
    .X(_08837_));
 sky130_fd_sc_hd__nand2_1 _15257_ (.A(_08837_),
    .B(_07848_),
    .Y(_08838_));
 sky130_fd_sc_hd__mux2_1 _15258_ (.A0(\core.cpuregs[24][21] ),
    .A1(\core.cpuregs[25][21] ),
    .S(_06240_),
    .X(_08839_));
 sky130_fd_sc_hd__mux2_1 _15259_ (.A0(\core.cpuregs[26][21] ),
    .A1(\core.cpuregs[27][21] ),
    .S(_06243_),
    .X(_08840_));
 sky130_fd_sc_hd__mux2_1 _15260_ (.A0(_08839_),
    .A1(_08840_),
    .S(_08253_),
    .X(_08841_));
 sky130_fd_sc_hd__mux2_1 _15261_ (.A0(\core.cpuregs[28][21] ),
    .A1(\core.cpuregs[29][21] ),
    .S(_06256_),
    .X(_08842_));
 sky130_fd_sc_hd__mux2_4 _15262_ (.A0(\core.cpuregs[30][21] ),
    .A1(\core.cpuregs[31][21] ),
    .S(_06250_),
    .X(_08843_));
 sky130_fd_sc_hd__mux2_1 _15263_ (.A0(_08842_),
    .A1(_08843_),
    .S(_06247_),
    .X(_08844_));
 sky130_fd_sc_hd__mux2_1 _15264_ (.A0(_08841_),
    .A1(_08844_),
    .S(_08249_),
    .X(_08845_));
 sky130_fd_sc_hd__mux2_1 _15265_ (.A0(\core.cpuregs[16][21] ),
    .A1(\core.cpuregs[17][21] ),
    .S(_06260_),
    .X(_08846_));
 sky130_fd_sc_hd__mux2_4 _15266_ (.A0(\core.cpuregs[18][21] ),
    .A1(\core.cpuregs[19][21] ),
    .S(_06273_),
    .X(_08847_));
 sky130_fd_sc_hd__mux2_1 _15267_ (.A0(_08846_),
    .A1(_08847_),
    .S(_06264_),
    .X(_08848_));
 sky130_fd_sc_hd__mux2_1 _15268_ (.A0(\core.cpuregs[22][21] ),
    .A1(\core.cpuregs[23][21] ),
    .S(_06273_),
    .X(_08849_));
 sky130_fd_sc_hd__mux2_1 _15269_ (.A0(\core.cpuregs[20][21] ),
    .A1(\core.cpuregs[21][21] ),
    .S(_06262_),
    .X(_08850_));
 sky130_fd_sc_hd__mux2_1 _15270_ (.A0(_08849_),
    .A1(_08850_),
    .S(_08257_),
    .X(_08851_));
 sky130_fd_sc_hd__mux2_8 _15271_ (.A0(_08848_),
    .A1(_08851_),
    .S(_06266_),
    .X(_08852_));
 sky130_fd_sc_hd__mux2_1 _15272_ (.A0(_08845_),
    .A1(_08852_),
    .S(_08558_),
    .X(_08853_));
 sky130_fd_sc_hd__nand2_1 _15273_ (.A(_08853_),
    .B(_07720_),
    .Y(_08854_));
 sky130_fd_sc_hd__a21o_1 _15274_ (.A1(_08838_),
    .A2(_08854_),
    .B1(_08561_),
    .X(_08855_));
 sky130_fd_sc_hd__or3b_1 _15275_ (.A(_08563_),
    .B(_08065_),
    .C_N(\core.reg_pc[21] ),
    .X(_08856_));
 sky130_fd_sc_hd__a21o_1 _15276_ (.A1(_08855_),
    .A2(_08856_),
    .B1(_07854_),
    .X(_08857_));
 sky130_fd_sc_hd__a21oi_1 _15277_ (.A1(_08814_),
    .A2(_06162_),
    .B1(_06159_),
    .Y(_08858_));
 sky130_fd_sc_hd__a31o_1 _15278_ (.A1(_08814_),
    .A2(_06159_),
    .A3(_06162_),
    .B1(_04395_),
    .X(_08859_));
 sky130_fd_sc_hd__or2_2 _15279_ (.A(_08858_),
    .B(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__nand2_1 _15280_ (.A(_08270_),
    .B(_04917_),
    .Y(_08861_));
 sky130_fd_sc_hd__and3_1 _15281_ (.A(_08861_),
    .B(_08571_),
    .C(_08714_),
    .X(_08862_));
 sky130_fd_sc_hd__nand2_1 _15282_ (.A(_08117_),
    .B(_04942_),
    .Y(_08863_));
 sky130_fd_sc_hd__and3_1 _15283_ (.A(_08272_),
    .B(_08712_),
    .C(_08863_),
    .X(_08864_));
 sky130_fd_sc_hd__o21ai_1 _15284_ (.A1(_08862_),
    .A2(_08864_),
    .B1(_08510_),
    .Y(_08865_));
 sky130_fd_sc_hd__nand3_1 _15285_ (.A(_08857_),
    .B(_08860_),
    .C(_08865_),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_1 _15286_ (.A(_08866_),
    .B(_08670_),
    .Y(_08867_));
 sky130_fd_sc_hd__o21ai_1 _15287_ (.A1(_04916_),
    .A2(_08773_),
    .B1(_08867_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand3_1 _15288_ (.A(_08812_),
    .B(_06160_),
    .C(_06163_),
    .Y(_08868_));
 sky130_fd_sc_hd__nand2_2 _15289_ (.A(_08868_),
    .B(_06186_),
    .Y(_08869_));
 sky130_fd_sc_hd__or2_1 _15290_ (.A(_06154_),
    .B(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__nand2_8 _15291_ (.A(_08869_),
    .B(_06154_),
    .Y(_08871_));
 sky130_fd_sc_hd__nand3_1 _15292_ (.A(_08870_),
    .B(_06225_),
    .C(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand2_1 _15293_ (.A(_07791_),
    .B(_04916_),
    .Y(_08873_));
 sky130_fd_sc_hd__and3_1 _15294_ (.A(_08873_),
    .B(_04626_),
    .C(_08764_),
    .X(_08874_));
 sky130_fd_sc_hd__nand2_1 _15295_ (.A(_07802_),
    .B(_04819_),
    .Y(_08875_));
 sky130_fd_sc_hd__and3_1 _15296_ (.A(_08272_),
    .B(_08762_),
    .C(_08875_),
    .X(_08876_));
 sky130_fd_sc_hd__o21ai_1 _15297_ (.A1(_08874_),
    .A2(_08876_),
    .B1(_05063_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand2_1 _15298_ (.A(_08872_),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__mux2_1 _15299_ (.A0(\core.cpuregs[12][22] ),
    .A1(\core.cpuregs[13][22] ),
    .S(_07773_),
    .X(_08879_));
 sky130_fd_sc_hd__clkbuf_2 _15300_ (.A(_07743_),
    .X(_08880_));
 sky130_fd_sc_hd__mux2_1 _15301_ (.A0(\core.cpuregs[14][22] ),
    .A1(\core.cpuregs[15][22] ),
    .S(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__mux2_1 _15302_ (.A0(_08879_),
    .A1(_08881_),
    .S(_07739_),
    .X(_08882_));
 sky130_fd_sc_hd__mux2_1 _15303_ (.A0(\core.cpuregs[8][22] ),
    .A1(\core.cpuregs[9][22] ),
    .S(_07773_),
    .X(_08883_));
 sky130_fd_sc_hd__mux2_2 _15304_ (.A0(\core.cpuregs[10][22] ),
    .A1(\core.cpuregs[11][22] ),
    .S(_08880_),
    .X(_08884_));
 sky130_fd_sc_hd__mux2_1 _15305_ (.A0(_08883_),
    .A1(_08884_),
    .S(_07739_),
    .X(_08885_));
 sky130_fd_sc_hd__mux2_1 _15306_ (.A0(_08882_),
    .A1(_08885_),
    .S(_07735_),
    .X(_08886_));
 sky130_fd_sc_hd__mux2_1 _15307_ (.A0(\core.cpuregs[0][22] ),
    .A1(\core.cpuregs[1][22] ),
    .S(_08880_),
    .X(_08887_));
 sky130_fd_sc_hd__mux2_2 _15308_ (.A0(\core.cpuregs[2][22] ),
    .A1(\core.cpuregs[3][22] ),
    .S(_07744_),
    .X(_08888_));
 sky130_fd_sc_hd__mux2_1 _15309_ (.A0(_08887_),
    .A1(_08888_),
    .S(_07664_),
    .X(_08889_));
 sky130_fd_sc_hd__mux2_1 _15310_ (.A0(\core.cpuregs[6][22] ),
    .A1(\core.cpuregs[7][22] ),
    .S(_07744_),
    .X(_08890_));
 sky130_fd_sc_hd__mux2_2 _15311_ (.A0(\core.cpuregs[4][22] ),
    .A1(\core.cpuregs[5][22] ),
    .S(_07744_),
    .X(_08891_));
 sky130_fd_sc_hd__mux2_1 _15312_ (.A0(_08890_),
    .A1(_08891_),
    .S(_07816_),
    .X(_08892_));
 sky130_fd_sc_hd__mux2_1 _15313_ (.A0(_08889_),
    .A1(_08892_),
    .S(_07741_),
    .X(_08893_));
 sky130_fd_sc_hd__mux2_1 _15314_ (.A0(_08886_),
    .A1(_08893_),
    .S(_07708_),
    .X(_08894_));
 sky130_fd_sc_hd__nand2_1 _15315_ (.A(_08894_),
    .B(_08739_),
    .Y(_08895_));
 sky130_fd_sc_hd__mux2_2 _15316_ (.A0(\core.cpuregs[24][22] ),
    .A1(\core.cpuregs[25][22] ),
    .S(_07746_),
    .X(_08896_));
 sky130_fd_sc_hd__clkbuf_2 _15317_ (.A(_07743_),
    .X(_08897_));
 sky130_fd_sc_hd__mux2_1 _15318_ (.A0(\core.cpuregs[26][22] ),
    .A1(\core.cpuregs[27][22] ),
    .S(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__mux2_1 _15319_ (.A0(_08896_),
    .A1(_08898_),
    .S(_07664_),
    .X(_08899_));
 sky130_fd_sc_hd__mux2_1 _15320_ (.A0(\core.cpuregs[28][22] ),
    .A1(\core.cpuregs[29][22] ),
    .S(_07746_),
    .X(_08900_));
 sky130_fd_sc_hd__mux2_1 _15321_ (.A0(\core.cpuregs[30][22] ),
    .A1(\core.cpuregs[31][22] ),
    .S(_08897_),
    .X(_08901_));
 sky130_fd_sc_hd__mux2_2 _15322_ (.A0(_08900_),
    .A1(_08901_),
    .S(_07754_),
    .X(_08902_));
 sky130_fd_sc_hd__mux2_8 _15323_ (.A0(_08899_),
    .A1(_08902_),
    .S(_07818_),
    .X(_08903_));
 sky130_fd_sc_hd__mux2_1 _15324_ (.A0(\core.cpuregs[16][22] ),
    .A1(\core.cpuregs[17][22] ),
    .S(_08897_),
    .X(_08904_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(\core.cpuregs[18][22] ),
    .A1(\core.cpuregs[19][22] ),
    .S(_07750_),
    .X(_08905_));
 sky130_fd_sc_hd__mux2_1 _15326_ (.A0(_08904_),
    .A1(_08905_),
    .S(_07754_),
    .X(_08906_));
 sky130_fd_sc_hd__mux2_1 _15327_ (.A0(\core.cpuregs[22][22] ),
    .A1(\core.cpuregs[23][22] ),
    .S(_07750_),
    .X(_08907_));
 sky130_fd_sc_hd__mux2_1 _15328_ (.A0(\core.cpuregs[20][22] ),
    .A1(\core.cpuregs[21][22] ),
    .S(_07750_),
    .X(_08908_));
 sky130_fd_sc_hd__mux2_1 _15329_ (.A0(_08907_),
    .A1(_08908_),
    .S(_07816_),
    .X(_08909_));
 sky130_fd_sc_hd__mux2_1 _15330_ (.A0(_08906_),
    .A1(_08909_),
    .S(_07818_),
    .X(_08910_));
 sky130_fd_sc_hd__mux2_1 _15331_ (.A0(_08903_),
    .A1(_08910_),
    .S(_07708_),
    .X(_08911_));
 sky130_fd_sc_hd__nand2_1 _15332_ (.A(_08911_),
    .B(_08756_),
    .Y(_08912_));
 sky130_fd_sc_hd__a21o_1 _15333_ (.A1(_08895_),
    .A2(_08912_),
    .B1(_07760_),
    .X(_08913_));
 sky130_fd_sc_hd__inv_2 _15334_ (.A(\core.reg_pc[22] ),
    .Y(_08914_));
 sky130_fd_sc_hd__or3_2 _15335_ (.A(_07729_),
    .B(_08914_),
    .C(_07852_),
    .X(_08915_));
 sky130_fd_sc_hd__a21oi_2 _15336_ (.A1(_08913_),
    .A2(_08915_),
    .B1(_08169_),
    .Y(_08916_));
 sky130_fd_sc_hd__o21ai_1 _15337_ (.A1(_08878_),
    .A2(_08916_),
    .B1(_07725_),
    .Y(_08917_));
 sky130_fd_sc_hd__o21ai_1 _15338_ (.A1(_04924_),
    .A2(_08773_),
    .B1(_08917_),
    .Y(_00265_));
 sky130_fd_sc_hd__mux2_1 _15339_ (.A0(\core.cpuregs[12][23] ),
    .A1(\core.cpuregs[13][23] ),
    .S(_08733_),
    .X(_08918_));
 sky130_fd_sc_hd__clkbuf_4 _15340_ (.A(_07691_),
    .X(_08919_));
 sky130_fd_sc_hd__mux2_1 _15341_ (.A0(\core.cpuregs[14][23] ),
    .A1(\core.cpuregs[15][23] ),
    .S(_08919_),
    .X(_08920_));
 sky130_fd_sc_hd__clkbuf_4 _15342_ (.A(_08285_),
    .X(_08921_));
 sky130_fd_sc_hd__mux2_1 _15343_ (.A0(_08918_),
    .A1(_08920_),
    .S(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__mux2_2 _15344_ (.A0(\core.cpuregs[8][23] ),
    .A1(\core.cpuregs[9][23] ),
    .S(_08733_),
    .X(_08923_));
 sky130_fd_sc_hd__clkbuf_4 _15345_ (.A(_07691_),
    .X(_08924_));
 sky130_fd_sc_hd__mux2_1 _15346_ (.A0(\core.cpuregs[10][23] ),
    .A1(\core.cpuregs[11][23] ),
    .S(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__mux2_1 _15347_ (.A0(_08923_),
    .A1(_08925_),
    .S(_08921_),
    .X(_08926_));
 sky130_fd_sc_hd__mux2_1 _15348_ (.A0(_08922_),
    .A1(_08926_),
    .S(_07696_),
    .X(_08927_));
 sky130_fd_sc_hd__mux2_1 _15349_ (.A0(\core.cpuregs[0][23] ),
    .A1(\core.cpuregs[1][23] ),
    .S(_08919_),
    .X(_08928_));
 sky130_fd_sc_hd__clkbuf_2 _15350_ (.A(_08514_),
    .X(_08929_));
 sky130_fd_sc_hd__mux2_1 _15351_ (.A0(\core.cpuregs[2][23] ),
    .A1(\core.cpuregs[3][23] ),
    .S(_08929_),
    .X(_08930_));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(_08928_),
    .A1(_08930_),
    .S(_08519_),
    .X(_08931_));
 sky130_fd_sc_hd__mux2_1 _15353_ (.A0(\core.cpuregs[6][23] ),
    .A1(\core.cpuregs[7][23] ),
    .S(_08924_),
    .X(_08932_));
 sky130_fd_sc_hd__mux2_1 _15354_ (.A0(\core.cpuregs[4][23] ),
    .A1(\core.cpuregs[5][23] ),
    .S(_08929_),
    .X(_08933_));
 sky130_fd_sc_hd__mux2_1 _15355_ (.A0(_08932_),
    .A1(_08933_),
    .S(_07694_),
    .X(_08934_));
 sky130_fd_sc_hd__mux2_1 _15356_ (.A0(_08931_),
    .A1(_08934_),
    .S(_08606_),
    .X(_08935_));
 sky130_fd_sc_hd__mux2_1 _15357_ (.A0(_08927_),
    .A1(_08935_),
    .S(_08737_),
    .X(_08936_));
 sky130_fd_sc_hd__nand2_1 _15358_ (.A(_08936_),
    .B(_08739_),
    .Y(_08937_));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(\core.cpuregs[24][23] ),
    .A1(\core.cpuregs[25][23] ),
    .S(_08649_),
    .X(_08938_));
 sky130_fd_sc_hd__clkbuf_4 _15360_ (.A(_08336_),
    .X(_08939_));
 sky130_fd_sc_hd__mux2_2 _15361_ (.A0(\core.cpuregs[26][23] ),
    .A1(\core.cpuregs[27][23] ),
    .S(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__clkbuf_4 _15362_ (.A(_06246_),
    .X(_08941_));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(_08938_),
    .A1(_08940_),
    .S(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__mux2_1 _15364_ (.A0(\core.cpuregs[28][23] ),
    .A1(\core.cpuregs[29][23] ),
    .S(_08939_),
    .X(_08943_));
 sky130_fd_sc_hd__buf_2 _15365_ (.A(_08336_),
    .X(_08944_));
 sky130_fd_sc_hd__mux2_1 _15366_ (.A0(\core.cpuregs[30][23] ),
    .A1(\core.cpuregs[31][23] ),
    .S(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(_08943_),
    .A1(_08945_),
    .S(_08941_),
    .X(_08946_));
 sky130_fd_sc_hd__mux2_1 _15368_ (.A0(_08942_),
    .A1(_08946_),
    .S(_08652_),
    .X(_08947_));
 sky130_fd_sc_hd__mux2_1 _15369_ (.A0(\core.cpuregs[16][23] ),
    .A1(\core.cpuregs[17][23] ),
    .S(_08944_),
    .X(_08948_));
 sky130_fd_sc_hd__clkbuf_4 _15370_ (.A(_08336_),
    .X(_08949_));
 sky130_fd_sc_hd__mux2_1 _15371_ (.A0(\core.cpuregs[18][23] ),
    .A1(\core.cpuregs[19][23] ),
    .S(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__mux2_1 _15372_ (.A0(_08948_),
    .A1(_08950_),
    .S(_08221_),
    .X(_08951_));
 sky130_fd_sc_hd__mux2_1 _15373_ (.A0(\core.cpuregs[22][23] ),
    .A1(\core.cpuregs[23][23] ),
    .S(_08949_),
    .X(_08952_));
 sky130_fd_sc_hd__mux2_1 _15374_ (.A0(\core.cpuregs[20][23] ),
    .A1(\core.cpuregs[21][23] ),
    .S(_08217_),
    .X(_08953_));
 sky130_fd_sc_hd__mux2_1 _15375_ (.A0(_08952_),
    .A1(_08953_),
    .S(_08247_),
    .X(_08954_));
 sky130_fd_sc_hd__mux2_2 _15376_ (.A0(_08951_),
    .A1(_08954_),
    .S(_08238_),
    .X(_08955_));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(_08947_),
    .A1(_08955_),
    .S(_08558_),
    .X(_08956_));
 sky130_fd_sc_hd__nand2_1 _15378_ (.A(_08956_),
    .B(_08756_),
    .Y(_08957_));
 sky130_fd_sc_hd__a21o_1 _15379_ (.A1(_08937_),
    .A2(_08957_),
    .B1(_08561_),
    .X(_08958_));
 sky130_fd_sc_hd__or3b_2 _15380_ (.A(_08563_),
    .B(_08065_),
    .C_N(\core.reg_pc[23] ),
    .X(_08959_));
 sky130_fd_sc_hd__a21o_1 _15381_ (.A1(_08958_),
    .A2(_08959_),
    .B1(_07894_),
    .X(_08960_));
 sky130_fd_sc_hd__nand2_1 _15382_ (.A(_08871_),
    .B(_06153_),
    .Y(_08961_));
 sky130_fd_sc_hd__or2_1 _15383_ (.A(_06151_),
    .B(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__nand2_1 _15384_ (.A(_08961_),
    .B(_06151_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand3_2 _15385_ (.A(_08962_),
    .B(_06226_),
    .C(_08963_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(_07790_),
    .B(_04924_),
    .Y(_08965_));
 sky130_fd_sc_hd__and3_1 _15387_ (.A(_08965_),
    .B(_08356_),
    .C(_08818_),
    .X(_08966_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_07787_),
    .B(_04814_),
    .Y(_08967_));
 sky130_fd_sc_hd__and3_1 _15389_ (.A(_07660_),
    .B(_08816_),
    .C(_08967_),
    .X(_08968_));
 sky130_fd_sc_hd__o21ai_1 _15390_ (.A1(_08966_),
    .A2(_08968_),
    .B1(_04634_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand3_1 _15391_ (.A(_08960_),
    .B(_08964_),
    .C(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__nand2_1 _15392_ (.A(_08970_),
    .B(_07725_),
    .Y(_08971_));
 sky130_fd_sc_hd__nand2_1 _15393_ (.A(_07728_),
    .B(_04879_),
    .Y(_08972_));
 sky130_fd_sc_hd__nand2_1 _15394_ (.A(_08971_),
    .B(_08972_),
    .Y(_00266_));
 sky130_fd_sc_hd__mux2_1 _15395_ (.A0(\core.cpuregs[12][24] ),
    .A1(\core.cpuregs[13][24] ),
    .S(_08288_),
    .X(_08973_));
 sky130_fd_sc_hd__mux2_1 _15396_ (.A0(\core.cpuregs[14][24] ),
    .A1(\core.cpuregs[15][24] ),
    .S(_08315_),
    .X(_08974_));
 sky130_fd_sc_hd__mux2_1 _15397_ (.A0(_08973_),
    .A1(_08974_),
    .S(_08302_),
    .X(_08975_));
 sky130_fd_sc_hd__mux2_1 _15398_ (.A0(\core.cpuregs[8][24] ),
    .A1(\core.cpuregs[9][24] ),
    .S(_08298_),
    .X(_08976_));
 sky130_fd_sc_hd__mux2_1 _15399_ (.A0(\core.cpuregs[10][24] ),
    .A1(\core.cpuregs[11][24] ),
    .S(_08300_),
    .X(_08977_));
 sky130_fd_sc_hd__mux2_1 _15400_ (.A0(_08976_),
    .A1(_08977_),
    .S(_08319_),
    .X(_08978_));
 sky130_fd_sc_hd__mux2_1 _15401_ (.A0(_08975_),
    .A1(_08978_),
    .S(_08417_),
    .X(_08979_));
 sky130_fd_sc_hd__mux2_1 _15402_ (.A0(\core.cpuregs[24][24] ),
    .A1(\core.cpuregs[25][24] ),
    .S(_08283_),
    .X(_08980_));
 sky130_fd_sc_hd__mux2_1 _15403_ (.A0(\core.cpuregs[26][24] ),
    .A1(\core.cpuregs[27][24] ),
    .S(_08329_),
    .X(_08981_));
 sky130_fd_sc_hd__mux2_4 _15404_ (.A0(_08980_),
    .A1(_08981_),
    .S(_08294_),
    .X(_08982_));
 sky130_fd_sc_hd__mux2_1 _15405_ (.A0(\core.cpuregs[28][24] ),
    .A1(\core.cpuregs[29][24] ),
    .S(_08422_),
    .X(_08983_));
 sky130_fd_sc_hd__mux2_1 _15406_ (.A0(\core.cpuregs[30][24] ),
    .A1(\core.cpuregs[31][24] ),
    .S(_08424_),
    .X(_08984_));
 sky130_fd_sc_hd__mux2_1 _15407_ (.A0(_08983_),
    .A1(_08984_),
    .S(_08332_),
    .X(_08985_));
 sky130_fd_sc_hd__mux2_1 _15408_ (.A0(_08982_),
    .A1(_08985_),
    .S(_08327_),
    .X(_08986_));
 sky130_fd_sc_hd__mux2_1 _15409_ (.A0(_08979_),
    .A1(_08986_),
    .S(_08343_),
    .X(_08987_));
 sky130_fd_sc_hd__mux2_2 _15410_ (.A0(\core.cpuregs[0][24] ),
    .A1(\core.cpuregs[1][24] ),
    .S(_08304_),
    .X(_08988_));
 sky130_fd_sc_hd__mux2_1 _15411_ (.A0(\core.cpuregs[2][24] ),
    .A1(\core.cpuregs[3][24] ),
    .S(_08307_),
    .X(_08989_));
 sky130_fd_sc_hd__mux2_1 _15412_ (.A0(_08988_),
    .A1(_08989_),
    .S(_08309_),
    .X(_08990_));
 sky130_fd_sc_hd__mux2_1 _15413_ (.A0(\core.cpuregs[6][24] ),
    .A1(\core.cpuregs[7][24] ),
    .S(_08317_),
    .X(_08991_));
 sky130_fd_sc_hd__mux2_1 _15414_ (.A0(\core.cpuregs[4][24] ),
    .A1(\core.cpuregs[5][24] ),
    .S(_08337_),
    .X(_08992_));
 sky130_fd_sc_hd__mux2_1 _15415_ (.A0(_08991_),
    .A1(_08992_),
    .S(_08339_),
    .X(_08993_));
 sky130_fd_sc_hd__mux2_1 _15416_ (.A0(_08990_),
    .A1(_08993_),
    .S(_08341_),
    .X(_08994_));
 sky130_fd_sc_hd__mux2_1 _15417_ (.A0(\core.cpuregs[16][24] ),
    .A1(\core.cpuregs[17][24] ),
    .S(_08321_),
    .X(_08995_));
 sky130_fd_sc_hd__mux2_1 _15418_ (.A0(\core.cpuregs[18][24] ),
    .A1(\core.cpuregs[19][24] ),
    .S(_08337_),
    .X(_08996_));
 sky130_fd_sc_hd__mux2_1 _15419_ (.A0(_08995_),
    .A1(_08996_),
    .S(_08438_),
    .X(_08997_));
 sky130_fd_sc_hd__mux2_1 _15420_ (.A0(\core.cpuregs[22][24] ),
    .A1(\core.cpuregs[23][24] ),
    .S(_08323_),
    .X(_08998_));
 sky130_fd_sc_hd__mux2_1 _15421_ (.A0(\core.cpuregs[20][24] ),
    .A1(\core.cpuregs[21][24] ),
    .S(_08649_),
    .X(_08999_));
 sky130_fd_sc_hd__mux2_1 _15422_ (.A0(_08998_),
    .A1(_08999_),
    .S(_08247_),
    .X(_09000_));
 sky130_fd_sc_hd__mux2_1 _15423_ (.A0(_08997_),
    .A1(_09000_),
    .S(_08652_),
    .X(_09001_));
 sky130_fd_sc_hd__mux2_1 _15424_ (.A0(_08994_),
    .A1(_09001_),
    .S(_08240_),
    .X(_09002_));
 sky130_fd_sc_hd__mux2_1 _15425_ (.A0(_08987_),
    .A1(_09002_),
    .S(_06293_),
    .X(_09003_));
 sky130_fd_sc_hd__nand2_1 _15426_ (.A(_09003_),
    .B(_07722_),
    .Y(_09004_));
 sky130_fd_sc_hd__inv_2 _15427_ (.A(\core.reg_pc[24] ),
    .Y(_09005_));
 sky130_fd_sc_hd__or3_1 _15428_ (.A(_06302_),
    .B(_09005_),
    .C(_06305_),
    .X(_09006_));
 sky130_fd_sc_hd__nand2_1 _15429_ (.A(_09004_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__nand2_1 _15430_ (.A(_09007_),
    .B(_06309_),
    .Y(_09008_));
 sky130_fd_sc_hd__or2_1 _15431_ (.A(_06202_),
    .B(_06189_),
    .X(_09009_));
 sky130_fd_sc_hd__nand2_8 _15432_ (.A(_06189_),
    .B(_06202_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand3_2 _15433_ (.A(_09009_),
    .B(_08503_),
    .C(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_1 _15434_ (.A(_08270_),
    .B(_04922_),
    .Y(_09012_));
 sky130_fd_sc_hd__and3_1 _15435_ (.A(_09012_),
    .B(_08571_),
    .C(_08863_),
    .X(_09013_));
 sky130_fd_sc_hd__nand2_1 _15436_ (.A(_08358_),
    .B(_04931_),
    .Y(_09014_));
 sky130_fd_sc_hd__and3_1 _15437_ (.A(_08272_),
    .B(_08861_),
    .C(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__o21ai_1 _15438_ (.A1(_09013_),
    .A2(_09015_),
    .B1(_05063_),
    .Y(_09016_));
 sky130_fd_sc_hd__nand3_1 _15439_ (.A(_09008_),
    .B(_09011_),
    .C(_09016_),
    .Y(_09017_));
 sky130_fd_sc_hd__nand2_1 _15440_ (.A(_09017_),
    .B(_08670_),
    .Y(_09018_));
 sky130_fd_sc_hd__o21ai_2 _15441_ (.A1(_04939_),
    .A2(_08773_),
    .B1(_09018_),
    .Y(_00267_));
 sky130_fd_sc_hd__mux2_1 _15442_ (.A0(\core.cpuregs[12][25] ),
    .A1(\core.cpuregs[13][25] ),
    .S(_07692_),
    .X(_09019_));
 sky130_fd_sc_hd__mux2_1 _15443_ (.A0(\core.cpuregs[14][25] ),
    .A1(\core.cpuregs[15][25] ),
    .S(_08720_),
    .X(_09020_));
 sky130_fd_sc_hd__mux2_1 _15444_ (.A0(_09019_),
    .A1(_09020_),
    .S(_08722_),
    .X(_09021_));
 sky130_fd_sc_hd__mux2_1 _15445_ (.A0(\core.cpuregs[8][25] ),
    .A1(\core.cpuregs[9][25] ),
    .S(_08720_),
    .X(_09022_));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(\core.cpuregs[10][25] ),
    .A1(\core.cpuregs[11][25] ),
    .S(_08725_),
    .X(_09023_));
 sky130_fd_sc_hd__mux2_1 _15447_ (.A0(_09022_),
    .A1(_09023_),
    .S(_08722_),
    .X(_09024_));
 sky130_fd_sc_hd__mux2_1 _15448_ (.A0(_09021_),
    .A1(_09024_),
    .S(_07696_),
    .X(_09025_));
 sky130_fd_sc_hd__mux2_1 _15449_ (.A0(\core.cpuregs[0][25] ),
    .A1(\core.cpuregs[1][25] ),
    .S(_08720_),
    .X(_09026_));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(\core.cpuregs[2][25] ),
    .A1(\core.cpuregs[3][25] ),
    .S(_08725_),
    .X(_09027_));
 sky130_fd_sc_hd__mux2_1 _15451_ (.A0(_09026_),
    .A1(_09027_),
    .S(_08722_),
    .X(_09028_));
 sky130_fd_sc_hd__mux2_1 _15452_ (.A0(\core.cpuregs[6][25] ),
    .A1(\core.cpuregs[7][25] ),
    .S(_08725_),
    .X(_09029_));
 sky130_fd_sc_hd__mux2_1 _15453_ (.A0(\core.cpuregs[4][25] ),
    .A1(\core.cpuregs[5][25] ),
    .S(_08733_),
    .X(_09030_));
 sky130_fd_sc_hd__mux2_1 _15454_ (.A0(_09029_),
    .A1(_09030_),
    .S(_07694_),
    .X(_09031_));
 sky130_fd_sc_hd__mux2_1 _15455_ (.A0(_09028_),
    .A1(_09031_),
    .S(_08606_),
    .X(_09032_));
 sky130_fd_sc_hd__mux2_1 _15456_ (.A0(_09025_),
    .A1(_09032_),
    .S(_08737_),
    .X(_09033_));
 sky130_fd_sc_hd__nand2_1 _15457_ (.A(_09033_),
    .B(_08739_),
    .Y(_09034_));
 sky130_fd_sc_hd__mux2_1 _15458_ (.A0(\core.cpuregs[24][25] ),
    .A1(\core.cpuregs[25][25] ),
    .S(_08517_),
    .X(_09035_));
 sky130_fd_sc_hd__mux2_1 _15459_ (.A0(\core.cpuregs[26][25] ),
    .A1(\core.cpuregs[27][25] ),
    .S(_08527_),
    .X(_09036_));
 sky130_fd_sc_hd__mux2_1 _15460_ (.A0(_09035_),
    .A1(_09036_),
    .S(_08524_),
    .X(_09037_));
 sky130_fd_sc_hd__mux2_1 _15461_ (.A0(\core.cpuregs[28][25] ),
    .A1(\core.cpuregs[29][25] ),
    .S(_08527_),
    .X(_09038_));
 sky130_fd_sc_hd__mux2_1 _15462_ (.A0(\core.cpuregs[30][25] ),
    .A1(\core.cpuregs[31][25] ),
    .S(_08533_),
    .X(_09039_));
 sky130_fd_sc_hd__mux2_2 _15463_ (.A0(_09038_),
    .A1(_09039_),
    .S(_08531_),
    .X(_09040_));
 sky130_fd_sc_hd__mux2_1 _15464_ (.A0(_09037_),
    .A1(_09040_),
    .S(_08539_),
    .X(_09041_));
 sky130_fd_sc_hd__mux2_1 _15465_ (.A0(\core.cpuregs[16][25] ),
    .A1(\core.cpuregs[17][25] ),
    .S(_08522_),
    .X(_09042_));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(\core.cpuregs[18][25] ),
    .A1(\core.cpuregs[19][25] ),
    .S(_08535_),
    .X(_09043_));
 sky130_fd_sc_hd__mux2_2 _15467_ (.A0(_09042_),
    .A1(_09043_),
    .S(_08531_),
    .X(_09044_));
 sky130_fd_sc_hd__mux2_1 _15468_ (.A0(\core.cpuregs[22][25] ),
    .A1(\core.cpuregs[23][25] ),
    .S(_08529_),
    .X(_09045_));
 sky130_fd_sc_hd__mux2_1 _15469_ (.A0(\core.cpuregs[20][25] ),
    .A1(\core.cpuregs[21][25] ),
    .S(_08535_),
    .X(_09046_));
 sky130_fd_sc_hd__mux2_2 _15470_ (.A0(_09045_),
    .A1(_09046_),
    .S(_08537_),
    .X(_09047_));
 sky130_fd_sc_hd__mux2_1 _15471_ (.A0(_09044_),
    .A1(_09047_),
    .S(_08311_),
    .X(_09048_));
 sky130_fd_sc_hd__mux2_1 _15472_ (.A0(_09041_),
    .A1(_09048_),
    .S(_08541_),
    .X(_09049_));
 sky130_fd_sc_hd__nand2_1 _15473_ (.A(_09049_),
    .B(_08756_),
    .Y(_09050_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(_09034_),
    .A2(_09050_),
    .B1(_07760_),
    .X(_09051_));
 sky130_fd_sc_hd__inv_2 _15475_ (.A(\core.reg_pc[25] ),
    .Y(_09052_));
 sky130_fd_sc_hd__or3_1 _15476_ (.A(_08563_),
    .B(_09052_),
    .C(_08496_),
    .X(_09053_));
 sky130_fd_sc_hd__nand2_1 _15477_ (.A(_09051_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _15478_ (.A(_07656_),
    .B(_04939_),
    .Y(_09055_));
 sky130_fd_sc_hd__and3_1 _15479_ (.A(_09055_),
    .B(_07902_),
    .C(_08875_),
    .X(_09056_));
 sky130_fd_sc_hd__nand2_1 _15480_ (.A(_07802_),
    .B(_04933_),
    .Y(_09057_));
 sky130_fd_sc_hd__and3_1 _15481_ (.A(_07786_),
    .B(_08873_),
    .C(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__o21a_1 _15482_ (.A1(_09056_),
    .A2(_09058_),
    .B1(_04633_),
    .X(_09059_));
 sky130_fd_sc_hd__a21oi_2 _15483_ (.A1(_09054_),
    .A2(_06309_),
    .B1(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_1 _15484_ (.A(_09010_),
    .B(_06201_),
    .Y(_09061_));
 sky130_fd_sc_hd__a21oi_1 _15485_ (.A1(_09061_),
    .A2(_06199_),
    .B1(_04984_),
    .Y(_09062_));
 sky130_fd_sc_hd__o21ai_2 _15486_ (.A1(_06199_),
    .A2(_09061_),
    .B1(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_8 _15487_ (.A(_09060_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__nand2_1 _15488_ (.A(_09064_),
    .B(_07652_),
    .Y(_09065_));
 sky130_fd_sc_hd__o21ai_2 _15489_ (.A1(_04942_),
    .A2(_08773_),
    .B1(_09065_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand3_1 _15490_ (.A(_06189_),
    .B(_06199_),
    .C(_06202_),
    .Y(_09066_));
 sky130_fd_sc_hd__nand2_1 _15491_ (.A(_09066_),
    .B(_06205_),
    .Y(_09067_));
 sky130_fd_sc_hd__or2_4 _15492_ (.A(_06193_),
    .B(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2_1 _15493_ (.A(_09067_),
    .B(_06193_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand3_1 _15494_ (.A(_09068_),
    .B(_06225_),
    .C(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_1 _15495_ (.A(_07790_),
    .B(_04942_),
    .Y(_09071_));
 sky130_fd_sc_hd__and3_1 _15496_ (.A(_09071_),
    .B(_04626_),
    .C(_08967_),
    .X(_09072_));
 sky130_fd_sc_hd__nand2_1 _15497_ (.A(_08117_),
    .B(_04843_),
    .Y(_09073_));
 sky130_fd_sc_hd__and3_1 _15498_ (.A(_07970_),
    .B(_08965_),
    .C(_09073_),
    .X(_09074_));
 sky130_fd_sc_hd__o21ai_1 _15499_ (.A1(_09072_),
    .A2(_09074_),
    .B1(_05063_),
    .Y(_09075_));
 sky130_fd_sc_hd__nand2_1 _15500_ (.A(_09070_),
    .B(_09075_),
    .Y(_09076_));
 sky130_fd_sc_hd__mux2_1 _15501_ (.A0(\core.cpuregs[12][26] ),
    .A1(\core.cpuregs[13][26] ),
    .S(_07773_),
    .X(_09077_));
 sky130_fd_sc_hd__mux2_1 _15502_ (.A0(\core.cpuregs[14][26] ),
    .A1(\core.cpuregs[15][26] ),
    .S(_08880_),
    .X(_09078_));
 sky130_fd_sc_hd__mux2_1 _15503_ (.A0(_09077_),
    .A1(_09078_),
    .S(_07739_),
    .X(_09079_));
 sky130_fd_sc_hd__mux2_1 _15504_ (.A0(\core.cpuregs[8][26] ),
    .A1(\core.cpuregs[9][26] ),
    .S(_07773_),
    .X(_09080_));
 sky130_fd_sc_hd__mux2_1 _15505_ (.A0(\core.cpuregs[10][26] ),
    .A1(\core.cpuregs[11][26] ),
    .S(_08880_),
    .X(_09081_));
 sky130_fd_sc_hd__mux2_1 _15506_ (.A0(_09080_),
    .A1(_09081_),
    .S(_07739_),
    .X(_09082_));
 sky130_fd_sc_hd__mux2_1 _15507_ (.A0(_09079_),
    .A1(_09082_),
    .S(_07735_),
    .X(_09083_));
 sky130_fd_sc_hd__mux2_1 _15508_ (.A0(\core.cpuregs[0][26] ),
    .A1(\core.cpuregs[1][26] ),
    .S(_08880_),
    .X(_09084_));
 sky130_fd_sc_hd__mux2_1 _15509_ (.A0(\core.cpuregs[2][26] ),
    .A1(\core.cpuregs[3][26] ),
    .S(_07744_),
    .X(_09085_));
 sky130_fd_sc_hd__mux2_1 _15510_ (.A0(_09084_),
    .A1(_09085_),
    .S(_07664_),
    .X(_09086_));
 sky130_fd_sc_hd__mux2_1 _15511_ (.A0(\core.cpuregs[6][26] ),
    .A1(\core.cpuregs[7][26] ),
    .S(_07744_),
    .X(_09087_));
 sky130_fd_sc_hd__mux2_1 _15512_ (.A0(\core.cpuregs[4][26] ),
    .A1(\core.cpuregs[5][26] ),
    .S(_07746_),
    .X(_09088_));
 sky130_fd_sc_hd__mux2_1 _15513_ (.A0(_09087_),
    .A1(_09088_),
    .S(_07816_),
    .X(_09089_));
 sky130_fd_sc_hd__mux2_1 _15514_ (.A0(_09086_),
    .A1(_09089_),
    .S(_07741_),
    .X(_09090_));
 sky130_fd_sc_hd__mux2_1 _15515_ (.A0(_09083_),
    .A1(_09090_),
    .S(_07708_),
    .X(_09091_));
 sky130_fd_sc_hd__nand2_1 _15516_ (.A(_09091_),
    .B(_08739_),
    .Y(_09092_));
 sky130_fd_sc_hd__mux2_1 _15517_ (.A0(\core.cpuregs[24][26] ),
    .A1(\core.cpuregs[25][26] ),
    .S(_07746_),
    .X(_09093_));
 sky130_fd_sc_hd__mux2_1 _15518_ (.A0(\core.cpuregs[26][26] ),
    .A1(\core.cpuregs[27][26] ),
    .S(_08897_),
    .X(_09094_));
 sky130_fd_sc_hd__mux2_4 _15519_ (.A0(_09093_),
    .A1(_09094_),
    .S(_07664_),
    .X(_09095_));
 sky130_fd_sc_hd__mux2_1 _15520_ (.A0(\core.cpuregs[28][26] ),
    .A1(\core.cpuregs[29][26] ),
    .S(_07746_),
    .X(_09096_));
 sky130_fd_sc_hd__mux2_1 _15521_ (.A0(\core.cpuregs[30][26] ),
    .A1(\core.cpuregs[31][26] ),
    .S(_08897_),
    .X(_09097_));
 sky130_fd_sc_hd__mux2_1 _15522_ (.A0(_09096_),
    .A1(_09097_),
    .S(_07754_),
    .X(_09098_));
 sky130_fd_sc_hd__mux2_1 _15523_ (.A0(_09095_),
    .A1(_09098_),
    .S(_07818_),
    .X(_09099_));
 sky130_fd_sc_hd__mux2_1 _15524_ (.A0(\core.cpuregs[16][26] ),
    .A1(\core.cpuregs[17][26] ),
    .S(_08897_),
    .X(_09100_));
 sky130_fd_sc_hd__mux2_1 _15525_ (.A0(\core.cpuregs[18][26] ),
    .A1(\core.cpuregs[19][26] ),
    .S(_07750_),
    .X(_09101_));
 sky130_fd_sc_hd__mux2_1 _15526_ (.A0(_09100_),
    .A1(_09101_),
    .S(_07754_),
    .X(_09102_));
 sky130_fd_sc_hd__mux2_1 _15527_ (.A0(\core.cpuregs[22][26] ),
    .A1(\core.cpuregs[23][26] ),
    .S(_07750_),
    .X(_09103_));
 sky130_fd_sc_hd__mux2_1 _15528_ (.A0(\core.cpuregs[20][26] ),
    .A1(\core.cpuregs[21][26] ),
    .S(_07752_),
    .X(_09104_));
 sky130_fd_sc_hd__mux2_1 _15529_ (.A0(_09103_),
    .A1(_09104_),
    .S(_07816_),
    .X(_09105_));
 sky130_fd_sc_hd__mux2_1 _15530_ (.A0(_09102_),
    .A1(_09105_),
    .S(_07818_),
    .X(_09106_));
 sky130_fd_sc_hd__mux2_1 _15531_ (.A0(_09099_),
    .A1(_09106_),
    .S(_07708_),
    .X(_09107_));
 sky130_fd_sc_hd__nand2_1 _15532_ (.A(_09107_),
    .B(_08756_),
    .Y(_09108_));
 sky130_fd_sc_hd__a21o_1 _15533_ (.A1(_09092_),
    .A2(_09108_),
    .B1(_07760_),
    .X(_09109_));
 sky130_fd_sc_hd__or3b_1 _15534_ (.A(_07729_),
    .B(_07852_),
    .C_N(_05464_),
    .X(_09110_));
 sky130_fd_sc_hd__a21oi_2 _15535_ (.A1(_09109_),
    .A2(_09110_),
    .B1(_08169_),
    .Y(_09111_));
 sky130_fd_sc_hd__o21ai_1 _15536_ (.A1(_09076_),
    .A2(_09111_),
    .B1(_07725_),
    .Y(_09112_));
 sky130_fd_sc_hd__o21ai_1 _15537_ (.A1(_04819_),
    .A2(_08773_),
    .B1(_09112_),
    .Y(_00269_));
 sky130_fd_sc_hd__mux2_1 _15538_ (.A0(\core.cpuregs[12][27] ),
    .A1(\core.cpuregs[13][27] ),
    .S(_08733_),
    .X(_09113_));
 sky130_fd_sc_hd__mux2_1 _15539_ (.A0(\core.cpuregs[14][27] ),
    .A1(\core.cpuregs[15][27] ),
    .S(_08919_),
    .X(_09114_));
 sky130_fd_sc_hd__mux2_1 _15540_ (.A0(_09113_),
    .A1(_09114_),
    .S(_08921_),
    .X(_09115_));
 sky130_fd_sc_hd__mux2_1 _15541_ (.A0(\core.cpuregs[8][27] ),
    .A1(\core.cpuregs[9][27] ),
    .S(_08919_),
    .X(_09116_));
 sky130_fd_sc_hd__mux2_4 _15542_ (.A0(\core.cpuregs[10][27] ),
    .A1(\core.cpuregs[11][27] ),
    .S(_08924_),
    .X(_09117_));
 sky130_fd_sc_hd__mux2_1 _15543_ (.A0(_09116_),
    .A1(_09117_),
    .S(_08921_),
    .X(_09118_));
 sky130_fd_sc_hd__mux2_1 _15544_ (.A0(_09115_),
    .A1(_09118_),
    .S(_08296_),
    .X(_09119_));
 sky130_fd_sc_hd__mux2_1 _15545_ (.A0(\core.cpuregs[0][27] ),
    .A1(\core.cpuregs[1][27] ),
    .S(_08924_),
    .X(_09120_));
 sky130_fd_sc_hd__mux2_2 _15546_ (.A0(\core.cpuregs[2][27] ),
    .A1(\core.cpuregs[3][27] ),
    .S(_08929_),
    .X(_09121_));
 sky130_fd_sc_hd__mux2_1 _15547_ (.A0(_09120_),
    .A1(_09121_),
    .S(_08519_),
    .X(_09122_));
 sky130_fd_sc_hd__mux2_1 _15548_ (.A0(\core.cpuregs[6][27] ),
    .A1(\core.cpuregs[7][27] ),
    .S(_08929_),
    .X(_09123_));
 sky130_fd_sc_hd__mux2_1 _15549_ (.A0(\core.cpuregs[4][27] ),
    .A1(\core.cpuregs[5][27] ),
    .S(_08515_),
    .X(_09124_));
 sky130_fd_sc_hd__mux2_1 _15550_ (.A0(_09123_),
    .A1(_09124_),
    .S(_07694_),
    .X(_09125_));
 sky130_fd_sc_hd__mux2_1 _15551_ (.A0(_09122_),
    .A1(_09125_),
    .S(_08606_),
    .X(_09126_));
 sky130_fd_sc_hd__mux2_1 _15552_ (.A0(_09119_),
    .A1(_09126_),
    .S(_08737_),
    .X(_09127_));
 sky130_fd_sc_hd__nand2_1 _15553_ (.A(_09127_),
    .B(_07848_),
    .Y(_09128_));
 sky130_fd_sc_hd__mux2_1 _15554_ (.A0(\core.cpuregs[24][27] ),
    .A1(\core.cpuregs[25][27] ),
    .S(_08649_),
    .X(_09129_));
 sky130_fd_sc_hd__mux2_1 _15555_ (.A0(\core.cpuregs[26][27] ),
    .A1(\core.cpuregs[27][27] ),
    .S(_08939_),
    .X(_09130_));
 sky130_fd_sc_hd__mux2_1 _15556_ (.A0(_09129_),
    .A1(_09130_),
    .S(_08941_),
    .X(_09131_));
 sky130_fd_sc_hd__mux2_2 _15557_ (.A0(\core.cpuregs[28][27] ),
    .A1(\core.cpuregs[29][27] ),
    .S(_08939_),
    .X(_09132_));
 sky130_fd_sc_hd__mux2_1 _15558_ (.A0(\core.cpuregs[30][27] ),
    .A1(\core.cpuregs[31][27] ),
    .S(_08944_),
    .X(_09133_));
 sky130_fd_sc_hd__mux2_1 _15559_ (.A0(_09132_),
    .A1(_09133_),
    .S(_08941_),
    .X(_09134_));
 sky130_fd_sc_hd__mux2_1 _15560_ (.A0(_09131_),
    .A1(_09134_),
    .S(_08652_),
    .X(_09135_));
 sky130_fd_sc_hd__mux2_1 _15561_ (.A0(\core.cpuregs[16][27] ),
    .A1(\core.cpuregs[17][27] ),
    .S(_08944_),
    .X(_09136_));
 sky130_fd_sc_hd__mux2_1 _15562_ (.A0(\core.cpuregs[18][27] ),
    .A1(\core.cpuregs[19][27] ),
    .S(_08949_),
    .X(_09137_));
 sky130_fd_sc_hd__mux2_1 _15563_ (.A0(_09136_),
    .A1(_09137_),
    .S(_08221_),
    .X(_09138_));
 sky130_fd_sc_hd__mux2_1 _15564_ (.A0(\core.cpuregs[22][27] ),
    .A1(\core.cpuregs[23][27] ),
    .S(_08949_),
    .X(_09139_));
 sky130_fd_sc_hd__mux2_1 _15565_ (.A0(\core.cpuregs[20][27] ),
    .A1(\core.cpuregs[21][27] ),
    .S(_08217_),
    .X(_09140_));
 sky130_fd_sc_hd__mux2_2 _15566_ (.A0(_09139_),
    .A1(_09140_),
    .S(_08247_),
    .X(_09141_));
 sky130_fd_sc_hd__mux2_1 _15567_ (.A0(_09138_),
    .A1(_09141_),
    .S(_08238_),
    .X(_09142_));
 sky130_fd_sc_hd__mux2_2 _15568_ (.A0(_09135_),
    .A1(_09142_),
    .S(_08558_),
    .X(_09143_));
 sky130_fd_sc_hd__nand2_8 _15569_ (.A(_09143_),
    .B(_07720_),
    .Y(_09144_));
 sky130_fd_sc_hd__a21o_1 _15570_ (.A1(_09128_),
    .A2(_09144_),
    .B1(_08561_),
    .X(_09145_));
 sky130_fd_sc_hd__or3b_2 _15571_ (.A(_08563_),
    .B(_08065_),
    .C_N(\core.reg_pc[27] ),
    .X(_09146_));
 sky130_fd_sc_hd__a21o_1 _15572_ (.A1(_09145_),
    .A2(_09146_),
    .B1(_07894_),
    .X(_09147_));
 sky130_fd_sc_hd__nand2_2 _15573_ (.A(_09069_),
    .B(_06192_),
    .Y(_09148_));
 sky130_fd_sc_hd__or2_1 _15574_ (.A(_06196_),
    .B(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__nand2_2 _15575_ (.A(_09148_),
    .B(_06196_),
    .Y(_09150_));
 sky130_fd_sc_hd__nand3_1 _15576_ (.A(_09149_),
    .B(_06226_),
    .C(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_1 _15577_ (.A(_07657_),
    .B(_04819_),
    .Y(_09152_));
 sky130_fd_sc_hd__and3_1 _15578_ (.A(_09152_),
    .B(_08356_),
    .C(_09014_),
    .X(_09153_));
 sky130_fd_sc_hd__nand2_1 _15579_ (.A(_06235_),
    .B(_04838_),
    .Y(_09154_));
 sky130_fd_sc_hd__and3_1 _15580_ (.A(_07660_),
    .B(_09012_),
    .C(_09154_),
    .X(_09155_));
 sky130_fd_sc_hd__o21ai_1 _15581_ (.A1(_09153_),
    .A2(_09155_),
    .B1(_04634_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand3_1 _15582_ (.A(_09147_),
    .B(_09151_),
    .C(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__nand2_1 _15583_ (.A(_09157_),
    .B(_07725_),
    .Y(_09158_));
 sky130_fd_sc_hd__nand2_2 _15584_ (.A(_07728_),
    .B(_06032_),
    .Y(_09159_));
 sky130_fd_sc_hd__nand2_1 _15585_ (.A(_09158_),
    .B(_09159_),
    .Y(_00270_));
 sky130_fd_sc_hd__mux2_1 _15586_ (.A0(\core.cpuregs[12][28] ),
    .A1(\core.cpuregs[13][28] ),
    .S(_07752_),
    .X(_09160_));
 sky130_fd_sc_hd__mux2_1 _15587_ (.A0(\core.cpuregs[14][28] ),
    .A1(\core.cpuregs[15][28] ),
    .S(_07752_),
    .X(_09161_));
 sky130_fd_sc_hd__mux2_1 _15588_ (.A0(_09160_),
    .A1(_09161_),
    .S(_07754_),
    .X(_09162_));
 sky130_fd_sc_hd__mux2_1 _15589_ (.A0(\core.cpuregs[8][28] ),
    .A1(\core.cpuregs[9][28] ),
    .S(_07752_),
    .X(_09163_));
 sky130_fd_sc_hd__mux2_1 _15590_ (.A0(\core.cpuregs[10][28] ),
    .A1(\core.cpuregs[11][28] ),
    .S(_07808_),
    .X(_09164_));
 sky130_fd_sc_hd__mux2_1 _15591_ (.A0(_09163_),
    .A1(_09164_),
    .S(_07812_),
    .X(_09165_));
 sky130_fd_sc_hd__mux2_1 _15592_ (.A0(_09162_),
    .A1(_09165_),
    .S(_07680_),
    .X(_09166_));
 sky130_fd_sc_hd__mux2_1 _15593_ (.A0(\core.cpuregs[0][28] ),
    .A1(\core.cpuregs[1][28] ),
    .S(_07752_),
    .X(_09167_));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(\core.cpuregs[2][28] ),
    .A1(\core.cpuregs[3][28] ),
    .S(_07808_),
    .X(_09168_));
 sky130_fd_sc_hd__mux2_1 _15595_ (.A0(_09167_),
    .A1(_09168_),
    .S(_07812_),
    .X(_09169_));
 sky130_fd_sc_hd__mux2_2 _15596_ (.A0(\core.cpuregs[6][28] ),
    .A1(\core.cpuregs[7][28] ),
    .S(_07808_),
    .X(_09170_));
 sky130_fd_sc_hd__mux2_2 _15597_ (.A0(\core.cpuregs[4][28] ),
    .A1(\core.cpuregs[5][28] ),
    .S(_07808_),
    .X(_09171_));
 sky130_fd_sc_hd__mux2_1 _15598_ (.A0(_09170_),
    .A1(_09171_),
    .S(_07816_),
    .X(_09172_));
 sky130_fd_sc_hd__mux2_1 _15599_ (.A0(_09169_),
    .A1(_09172_),
    .S(_07818_),
    .X(_09173_));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(_09166_),
    .A1(_09173_),
    .S(_08737_),
    .X(_09174_));
 sky130_fd_sc_hd__nand2_2 _15601_ (.A(_09174_),
    .B(_08739_),
    .Y(_09175_));
 sky130_fd_sc_hd__mux2_1 _15602_ (.A0(\core.cpuregs[24][28] ),
    .A1(\core.cpuregs[25][28] ),
    .S(_07835_),
    .X(_09176_));
 sky130_fd_sc_hd__mux2_1 _15603_ (.A0(\core.cpuregs[26][28] ),
    .A1(\core.cpuregs[27][28] ),
    .S(_07835_),
    .X(_09177_));
 sky130_fd_sc_hd__mux2_4 _15604_ (.A0(_09176_),
    .A1(_09177_),
    .S(_07841_),
    .X(_09178_));
 sky130_fd_sc_hd__mux2_2 _15605_ (.A0(\core.cpuregs[28][28] ),
    .A1(\core.cpuregs[29][28] ),
    .S(_07835_),
    .X(_09179_));
 sky130_fd_sc_hd__mux2_4 _15606_ (.A0(\core.cpuregs[30][28] ),
    .A1(\core.cpuregs[31][28] ),
    .S(_07906_),
    .X(_09180_));
 sky130_fd_sc_hd__mux2_1 _15607_ (.A0(_09179_),
    .A1(_09180_),
    .S(_07841_),
    .X(_09181_));
 sky130_fd_sc_hd__mux2_1 _15608_ (.A0(_09178_),
    .A1(_09181_),
    .S(_07828_),
    .X(_09182_));
 sky130_fd_sc_hd__mux2_1 _15609_ (.A0(\core.cpuregs[16][28] ),
    .A1(\core.cpuregs[17][28] ),
    .S(_07835_),
    .X(_09183_));
 sky130_fd_sc_hd__mux2_2 _15610_ (.A0(\core.cpuregs[18][28] ),
    .A1(\core.cpuregs[19][28] ),
    .S(_07906_),
    .X(_09184_));
 sky130_fd_sc_hd__mux2_1 _15611_ (.A0(_09183_),
    .A1(_09184_),
    .S(_07841_),
    .X(_09185_));
 sky130_fd_sc_hd__mux2_1 _15612_ (.A0(\core.cpuregs[22][28] ),
    .A1(\core.cpuregs[23][28] ),
    .S(_07906_),
    .X(_09186_));
 sky130_fd_sc_hd__mux2_1 _15613_ (.A0(\core.cpuregs[20][28] ),
    .A1(\core.cpuregs[21][28] ),
    .S(_07906_),
    .X(_09187_));
 sky130_fd_sc_hd__mux2_1 _15614_ (.A0(_09186_),
    .A1(_09187_),
    .S(_07671_),
    .X(_09188_));
 sky130_fd_sc_hd__mux2_1 _15615_ (.A0(_09185_),
    .A1(_09188_),
    .S(_07828_),
    .X(_09189_));
 sky130_fd_sc_hd__mux2_1 _15616_ (.A0(_09182_),
    .A1(_09189_),
    .S(_08737_),
    .X(_09190_));
 sky130_fd_sc_hd__nand2_1 _15617_ (.A(_09190_),
    .B(_08756_),
    .Y(_09191_));
 sky130_fd_sc_hd__a21o_1 _15618_ (.A1(_09175_),
    .A2(_09191_),
    .B1(_07760_),
    .X(_09192_));
 sky130_fd_sc_hd__inv_2 _15619_ (.A(_05492_),
    .Y(_09193_));
 sky130_fd_sc_hd__or3_1 _15620_ (.A(_07729_),
    .B(_09193_),
    .C(_07852_),
    .X(_09194_));
 sky130_fd_sc_hd__a21oi_1 _15621_ (.A1(_09192_),
    .A2(_09194_),
    .B1(_08169_),
    .Y(_09195_));
 sky130_fd_sc_hd__or2_1 _15622_ (.A(_06214_),
    .B(_06208_),
    .X(_09196_));
 sky130_fd_sc_hd__nand2_1 _15623_ (.A(_06208_),
    .B(_06214_),
    .Y(_09197_));
 sky130_fd_sc_hd__o211a_1 _15624_ (.A1(_06032_),
    .A2(_07802_),
    .B1(_09057_),
    .C1(_07902_),
    .X(_09198_));
 sky130_fd_sc_hd__o21ai_2 _15625_ (.A1(_04838_),
    .A2(_06231_),
    .B1(_06234_),
    .Y(_09199_));
 sky130_fd_sc_hd__and3_1 _15626_ (.A(_07659_),
    .B(_09055_),
    .C(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__o21a_1 _15627_ (.A1(_09198_),
    .A2(_09200_),
    .B1(_05062_),
    .X(_09201_));
 sky130_fd_sc_hd__a31o_1 _15628_ (.A1(_09196_),
    .A2(_06225_),
    .A3(_09197_),
    .B1(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__o21ai_1 _15629_ (.A1(_09195_),
    .A2(_09202_),
    .B1(_07980_),
    .Y(_09203_));
 sky130_fd_sc_hd__o21ai_1 _15630_ (.A1(_04931_),
    .A2(_07724_),
    .B1(_09203_),
    .Y(_00271_));
 sky130_fd_sc_hd__mux2_1 _15631_ (.A0(\core.cpuregs[12][29] ),
    .A1(\core.cpuregs[13][29] ),
    .S(_08515_),
    .X(_09204_));
 sky130_fd_sc_hd__mux2_1 _15632_ (.A0(\core.cpuregs[14][29] ),
    .A1(\core.cpuregs[15][29] ),
    .S(_08527_),
    .X(_09205_));
 sky130_fd_sc_hd__mux2_1 _15633_ (.A0(_09204_),
    .A1(_09205_),
    .S(_08519_),
    .X(_09206_));
 sky130_fd_sc_hd__mux2_1 _15634_ (.A0(\core.cpuregs[8][29] ),
    .A1(\core.cpuregs[9][29] ),
    .S(_08517_),
    .X(_09207_));
 sky130_fd_sc_hd__mux2_1 _15635_ (.A0(\core.cpuregs[10][29] ),
    .A1(\core.cpuregs[11][29] ),
    .S(_08533_),
    .X(_09208_));
 sky130_fd_sc_hd__mux2_1 _15636_ (.A0(_09207_),
    .A1(_09208_),
    .S(_08524_),
    .X(_09209_));
 sky130_fd_sc_hd__mux2_1 _15637_ (.A0(_09206_),
    .A1(_09209_),
    .S(_08296_),
    .X(_09210_));
 sky130_fd_sc_hd__mux2_1 _15638_ (.A0(\core.cpuregs[0][29] ),
    .A1(\core.cpuregs[1][29] ),
    .S(_08522_),
    .X(_09211_));
 sky130_fd_sc_hd__mux2_1 _15639_ (.A0(\core.cpuregs[2][29] ),
    .A1(\core.cpuregs[3][29] ),
    .S(_08529_),
    .X(_09212_));
 sky130_fd_sc_hd__mux2_1 _15640_ (.A0(_09211_),
    .A1(_09212_),
    .S(_08531_),
    .X(_09213_));
 sky130_fd_sc_hd__mux2_1 _15641_ (.A0(\core.cpuregs[6][29] ),
    .A1(\core.cpuregs[7][29] ),
    .S(_08533_),
    .X(_09214_));
 sky130_fd_sc_hd__mux2_2 _15642_ (.A0(\core.cpuregs[4][29] ),
    .A1(\core.cpuregs[5][29] ),
    .S(_08535_),
    .X(_09215_));
 sky130_fd_sc_hd__mux2_1 _15643_ (.A0(_09214_),
    .A1(_09215_),
    .S(_08537_),
    .X(_09216_));
 sky130_fd_sc_hd__mux2_1 _15644_ (.A0(_09213_),
    .A1(_09216_),
    .S(_08539_),
    .X(_09217_));
 sky130_fd_sc_hd__mux2_1 _15645_ (.A0(_09210_),
    .A1(_09217_),
    .S(_08541_),
    .X(_09218_));
 sky130_fd_sc_hd__nand2_1 _15646_ (.A(_09218_),
    .B(_07848_),
    .Y(_09219_));
 sky130_fd_sc_hd__mux2_1 _15647_ (.A0(\core.cpuregs[24][29] ),
    .A1(\core.cpuregs[25][29] ),
    .S(_06240_),
    .X(_09220_));
 sky130_fd_sc_hd__mux2_4 _15648_ (.A0(\core.cpuregs[26][29] ),
    .A1(\core.cpuregs[27][29] ),
    .S(_06243_),
    .X(_09221_));
 sky130_fd_sc_hd__mux2_1 _15649_ (.A0(_09220_),
    .A1(_09221_),
    .S(_08253_),
    .X(_09222_));
 sky130_fd_sc_hd__mux2_1 _15650_ (.A0(\core.cpuregs[28][29] ),
    .A1(\core.cpuregs[29][29] ),
    .S(_06256_),
    .X(_09223_));
 sky130_fd_sc_hd__mux2_1 _15651_ (.A0(\core.cpuregs[30][29] ),
    .A1(\core.cpuregs[31][29] ),
    .S(_06250_),
    .X(_09224_));
 sky130_fd_sc_hd__mux2_1 _15652_ (.A0(_09223_),
    .A1(_09224_),
    .S(_06247_),
    .X(_09225_));
 sky130_fd_sc_hd__mux2_1 _15653_ (.A0(_09222_),
    .A1(_09225_),
    .S(_06266_),
    .X(_09226_));
 sky130_fd_sc_hd__mux2_1 _15654_ (.A0(\core.cpuregs[16][29] ),
    .A1(\core.cpuregs[17][29] ),
    .S(_06260_),
    .X(_09227_));
 sky130_fd_sc_hd__mux2_2 _15655_ (.A0(\core.cpuregs[18][29] ),
    .A1(\core.cpuregs[19][29] ),
    .S(_06262_),
    .X(_09228_));
 sky130_fd_sc_hd__mux2_1 _15656_ (.A0(_09227_),
    .A1(_09228_),
    .S(_06264_),
    .X(_09229_));
 sky130_fd_sc_hd__mux2_1 _15657_ (.A0(\core.cpuregs[22][29] ),
    .A1(\core.cpuregs[23][29] ),
    .S(_06273_),
    .X(_09230_));
 sky130_fd_sc_hd__mux2_1 _15658_ (.A0(\core.cpuregs[20][29] ),
    .A1(\core.cpuregs[21][29] ),
    .S(_06276_),
    .X(_09231_));
 sky130_fd_sc_hd__mux2_1 _15659_ (.A0(_09230_),
    .A1(_09231_),
    .S(_08257_),
    .X(_09232_));
 sky130_fd_sc_hd__mux2_1 _15660_ (.A0(_09229_),
    .A1(_09232_),
    .S(_06266_),
    .X(_09233_));
 sky130_fd_sc_hd__mux2_1 _15661_ (.A0(_09226_),
    .A1(_09233_),
    .S(_08558_),
    .X(_09234_));
 sky130_fd_sc_hd__nand2_1 _15662_ (.A(_09234_),
    .B(_07720_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21o_1 _15663_ (.A1(_09219_),
    .A2(_09235_),
    .B1(_08561_),
    .X(_09236_));
 sky130_fd_sc_hd__inv_2 _15664_ (.A(\core.reg_pc[29] ),
    .Y(_09237_));
 sky130_fd_sc_hd__or3_1 _15665_ (.A(_07964_),
    .B(_09237_),
    .C(_08496_),
    .X(_09238_));
 sky130_fd_sc_hd__a21o_1 _15666_ (.A1(_09236_),
    .A2(_09238_),
    .B1(_07854_),
    .X(_09239_));
 sky130_fd_sc_hd__nand2_1 _15667_ (.A(_09197_),
    .B(_06213_),
    .Y(_09240_));
 sky130_fd_sc_hd__or2_1 _15668_ (.A(_06211_),
    .B(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__nand2_1 _15669_ (.A(_09240_),
    .B(_06211_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand3_1 _15670_ (.A(_09241_),
    .B(_08503_),
    .C(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__o211a_1 _15671_ (.A1(_04849_),
    .A2(_06235_),
    .B1(_09073_),
    .C1(_04589_),
    .X(_09244_));
 sky130_fd_sc_hd__and3_1 _15672_ (.A(_08272_),
    .B(_09071_),
    .C(_09199_),
    .X(_09245_));
 sky130_fd_sc_hd__o21ai_1 _15673_ (.A1(_09244_),
    .A2(_09245_),
    .B1(_05063_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand3_1 _15674_ (.A(_09239_),
    .B(_09243_),
    .C(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__nand2_1 _15675_ (.A(_09247_),
    .B(_07652_),
    .Y(_09248_));
 sky130_fd_sc_hd__o21ai_2 _15676_ (.A1(_04933_),
    .A2(_07724_),
    .B1(_09248_),
    .Y(_00272_));
 sky130_fd_sc_hd__mux2_1 _15677_ (.A0(\core.cpuregs[12][30] ),
    .A1(\core.cpuregs[13][30] ),
    .S(_08733_),
    .X(_09249_));
 sky130_fd_sc_hd__mux2_1 _15678_ (.A0(\core.cpuregs[14][30] ),
    .A1(\core.cpuregs[15][30] ),
    .S(_08919_),
    .X(_09250_));
 sky130_fd_sc_hd__mux2_1 _15679_ (.A0(_09249_),
    .A1(_09250_),
    .S(_08921_),
    .X(_09251_));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(\core.cpuregs[8][30] ),
    .A1(\core.cpuregs[9][30] ),
    .S(_08919_),
    .X(_09252_));
 sky130_fd_sc_hd__mux2_1 _15681_ (.A0(\core.cpuregs[10][30] ),
    .A1(\core.cpuregs[11][30] ),
    .S(_08924_),
    .X(_09253_));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(_09252_),
    .A1(_09253_),
    .S(_08921_),
    .X(_09254_));
 sky130_fd_sc_hd__mux2_1 _15683_ (.A0(_09251_),
    .A1(_09254_),
    .S(_08296_),
    .X(_09255_));
 sky130_fd_sc_hd__mux2_1 _15684_ (.A0(\core.cpuregs[0][30] ),
    .A1(\core.cpuregs[1][30] ),
    .S(_08924_),
    .X(_09256_));
 sky130_fd_sc_hd__mux2_1 _15685_ (.A0(\core.cpuregs[2][30] ),
    .A1(\core.cpuregs[3][30] ),
    .S(_08929_),
    .X(_09257_));
 sky130_fd_sc_hd__mux2_1 _15686_ (.A0(_09256_),
    .A1(_09257_),
    .S(_08519_),
    .X(_09258_));
 sky130_fd_sc_hd__mux2_1 _15687_ (.A0(\core.cpuregs[6][30] ),
    .A1(\core.cpuregs[7][30] ),
    .S(_08929_),
    .X(_09259_));
 sky130_fd_sc_hd__mux2_1 _15688_ (.A0(\core.cpuregs[4][30] ),
    .A1(\core.cpuregs[5][30] ),
    .S(_08515_),
    .X(_09260_));
 sky130_fd_sc_hd__mux2_1 _15689_ (.A0(_09259_),
    .A1(_09260_),
    .S(_08537_),
    .X(_09261_));
 sky130_fd_sc_hd__mux2_1 _15690_ (.A0(_09258_),
    .A1(_09261_),
    .S(_08606_),
    .X(_09262_));
 sky130_fd_sc_hd__mux2_1 _15691_ (.A0(_09255_),
    .A1(_09262_),
    .S(_08541_),
    .X(_09263_));
 sky130_fd_sc_hd__nand2_1 _15692_ (.A(_09263_),
    .B(_07848_),
    .Y(_09264_));
 sky130_fd_sc_hd__mux2_1 _15693_ (.A0(\core.cpuregs[24][30] ),
    .A1(\core.cpuregs[25][30] ),
    .S(_08939_),
    .X(_09265_));
 sky130_fd_sc_hd__mux2_1 _15694_ (.A0(\core.cpuregs[26][30] ),
    .A1(\core.cpuregs[27][30] ),
    .S(_08944_),
    .X(_09266_));
 sky130_fd_sc_hd__mux2_1 _15695_ (.A0(_09265_),
    .A1(_09266_),
    .S(_08941_),
    .X(_09267_));
 sky130_fd_sc_hd__mux2_1 _15696_ (.A0(\core.cpuregs[28][30] ),
    .A1(\core.cpuregs[29][30] ),
    .S(_08939_),
    .X(_09268_));
 sky130_fd_sc_hd__mux2_1 _15697_ (.A0(\core.cpuregs[30][30] ),
    .A1(\core.cpuregs[31][30] ),
    .S(_08949_),
    .X(_09269_));
 sky130_fd_sc_hd__mux2_1 _15698_ (.A0(_09268_),
    .A1(_09269_),
    .S(_08941_),
    .X(_09270_));
 sky130_fd_sc_hd__mux2_1 _15699_ (.A0(_09267_),
    .A1(_09270_),
    .S(_08238_),
    .X(_09271_));
 sky130_fd_sc_hd__mux2_1 _15700_ (.A0(\core.cpuregs[16][30] ),
    .A1(\core.cpuregs[17][30] ),
    .S(_08944_),
    .X(_09272_));
 sky130_fd_sc_hd__mux2_1 _15701_ (.A0(\core.cpuregs[18][30] ),
    .A1(\core.cpuregs[19][30] ),
    .S(_08217_),
    .X(_09273_));
 sky130_fd_sc_hd__mux2_1 _15702_ (.A0(_09272_),
    .A1(_09273_),
    .S(_08221_),
    .X(_09274_));
 sky130_fd_sc_hd__mux2_1 _15703_ (.A0(\core.cpuregs[22][30] ),
    .A1(\core.cpuregs[23][30] ),
    .S(_08949_),
    .X(_09275_));
 sky130_fd_sc_hd__mux2_1 _15704_ (.A0(\core.cpuregs[20][30] ),
    .A1(\core.cpuregs[21][30] ),
    .S(_08217_),
    .X(_09276_));
 sky130_fd_sc_hd__mux2_1 _15705_ (.A0(_09275_),
    .A1(_09276_),
    .S(_08247_),
    .X(_09277_));
 sky130_fd_sc_hd__mux2_1 _15706_ (.A0(_09274_),
    .A1(_09277_),
    .S(_08238_),
    .X(_09278_));
 sky130_fd_sc_hd__mux2_1 _15707_ (.A0(_09271_),
    .A1(_09278_),
    .S(_08558_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2_4 _15708_ (.A(_09279_),
    .B(_07720_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21o_1 _15709_ (.A1(_09264_),
    .A2(_09280_),
    .B1(_08561_),
    .X(_09281_));
 sky130_fd_sc_hd__or3_2 _15710_ (.A(_08563_),
    .B(_05518_),
    .C(_08496_),
    .X(_09282_));
 sky130_fd_sc_hd__a21o_1 _15711_ (.A1(_09281_),
    .A2(_09282_),
    .B1(_07894_),
    .X(_09283_));
 sky130_fd_sc_hd__or2_1 _15712_ (.A(_06220_),
    .B(_06217_),
    .X(_09284_));
 sky130_fd_sc_hd__nand3_1 _15713_ (.A(_09284_),
    .B(_06226_),
    .C(_06221_),
    .Y(_09285_));
 sky130_fd_sc_hd__o211a_1 _15714_ (.A1(_04856_),
    .A2(_06235_),
    .B1(_09154_),
    .C1(_04589_),
    .X(_09286_));
 sky130_fd_sc_hd__and3_1 _15715_ (.A(_07660_),
    .B(_09152_),
    .C(_09199_),
    .X(_09287_));
 sky130_fd_sc_hd__o21ai_1 _15716_ (.A1(_09286_),
    .A2(_09287_),
    .B1(_04634_),
    .Y(_09288_));
 sky130_fd_sc_hd__nand3_1 _15717_ (.A(_09283_),
    .B(_09285_),
    .C(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_2 _15718_ (.A(_09289_),
    .B(_07725_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_2 _15719_ (.A(_07728_),
    .B(_04845_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand2_8 _15720_ (.A(_09290_),
    .B(_09291_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _15721_ (.A(_04374_),
    .B(\core.mem_state[0] ),
    .Y(_09292_));
 sky130_fd_sc_hd__or3_1 _15722_ (.A(\core.mem_do_rinst ),
    .B(\core.mem_do_rdata ),
    .C(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_04371_),
    .B(_04370_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor2_1 _15724_ (.A(net103),
    .B(_04512_),
    .Y(_09295_));
 sky130_fd_sc_hd__inv_2 _15725_ (.A(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__buf_2 _15726_ (.A(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__a21oi_1 _15727_ (.A1(_09293_),
    .A2(_09294_),
    .B1(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__nand2_1 _15728_ (.A(_04375_),
    .B(\core.mem_state[1] ),
    .Y(_09299_));
 sky130_fd_sc_hd__a221o_1 _15729_ (.A1(net66),
    .A2(net33),
    .B1(_09292_),
    .B2(_09299_),
    .C1(_09297_),
    .X(_09300_));
 sky130_fd_sc_hd__o41a_2 _15730_ (.A1(\core.mem_do_rdata ),
    .A2(_05960_),
    .A3(_09297_),
    .A4(_09294_),
    .B1(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__nand2_2 _15731_ (.A(_04388_),
    .B(net103),
    .Y(_09302_));
 sky130_fd_sc_hd__or4_1 _15732_ (.A(\core.mem_do_rinst ),
    .B(_04374_),
    .C(_04375_),
    .D(_09297_),
    .X(_09303_));
 sky130_fd_sc_hd__nand3_2 _15733_ (.A(_09301_),
    .B(_09302_),
    .C(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__mux2_1 _15734_ (.A0(_09298_),
    .A1(\core.mem_state[0] ),
    .S(_09304_),
    .X(_09305_));
 sky130_fd_sc_hd__clkbuf_1 _15735_ (.A(_09305_),
    .X(_00274_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(_04371_),
    .B(\core.mem_do_wdata ),
    .Y(_09306_));
 sky130_fd_sc_hd__a21oi_1 _15737_ (.A1(_09293_),
    .A2(_09306_),
    .B1(_09297_),
    .Y(_09307_));
 sky130_fd_sc_hd__mux2_1 _15738_ (.A0(_09307_),
    .A1(\core.mem_state[1] ),
    .S(_09304_),
    .X(_09308_));
 sky130_fd_sc_hd__clkbuf_1 _15739_ (.A(_09308_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _15740_ (.A0(\core.reg_out[0] ),
    .A1(\core.alu_out_q[0] ),
    .S(_06601_),
    .X(_09309_));
 sky130_fd_sc_hd__inv_2 _15741_ (.A(\core.latched_store ),
    .Y(_09310_));
 sky130_fd_sc_hd__nor2_1 _15742_ (.A(\core.latched_branch ),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15743_ (.A(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15744_ (.A(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__and2_1 _15745_ (.A(_09309_),
    .B(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15746_ (.A(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__inv_2 _15747_ (.A(\core.latched_branch ),
    .Y(_09316_));
 sky130_fd_sc_hd__inv_2 _15748_ (.A(\core.latched_rd[4] ),
    .Y(_09317_));
 sky130_fd_sc_hd__inv_2 _15749_ (.A(\core.latched_rd[3] ),
    .Y(_09318_));
 sky130_fd_sc_hd__inv_2 _15750_ (.A(\core.latched_rd[2] ),
    .Y(_09319_));
 sky130_fd_sc_hd__and3_1 _15751_ (.A(_09317_),
    .B(_09318_),
    .C(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(\core.latched_rd[1] ),
    .B(\core.latched_rd[0] ),
    .Y(_09321_));
 sky130_fd_sc_hd__a221o_1 _15753_ (.A1(_09310_),
    .A2(_09316_),
    .B1(_09320_),
    .B2(_09321_),
    .C1(_04457_),
    .X(_09322_));
 sky130_fd_sc_hd__inv_2 _15754_ (.A(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__buf_1 _15755_ (.A(_09323_),
    .X(_09324_));
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(\core.latched_rd[1] ),
    .B(\core.latched_rd[0] ),
    .Y(_09325_));
 sky130_fd_sc_hd__inv_2 _15757_ (.A(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__or3_1 _15758_ (.A(\core.latched_rd[3] ),
    .B(_09317_),
    .C(_09319_),
    .X(_09327_));
 sky130_fd_sc_hd__inv_2 _15759_ (.A(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__and3_1 _15760_ (.A(_09324_),
    .B(_09326_),
    .C(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__buf_4 _15761_ (.A(_09329_),
    .X(_09330_));
 sky130_fd_sc_hd__clkbuf_4 _15762_ (.A(_09330_),
    .X(_09331_));
 sky130_fd_sc_hd__mux2_2 _15763_ (.A0(\core.cpuregs[23][0] ),
    .A1(_09315_),
    .S(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__buf_1 _15764_ (.A(_09332_),
    .X(_00276_));
 sky130_fd_sc_hd__nand2_1 _15765_ (.A(_06598_),
    .B(_06602_),
    .Y(_09333_));
 sky130_fd_sc_hd__buf_1 _15766_ (.A(_09311_),
    .X(_09334_));
 sky130_fd_sc_hd__clkbuf_2 _15767_ (.A(_09334_),
    .X(_09335_));
 sky130_fd_sc_hd__mux2_1 _15768_ (.A0(\core.reg_pc[1] ),
    .A1(_09333_),
    .S(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__buf_1 _15769_ (.A(_09336_),
    .X(_09337_));
 sky130_fd_sc_hd__mux2_1 _15770_ (.A0(\core.cpuregs[23][1] ),
    .A1(_09337_),
    .S(_09331_),
    .X(_09338_));
 sky130_fd_sc_hd__clkbuf_1 _15771_ (.A(_09338_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _15772_ (.A0(_05053_),
    .A1(_06622_),
    .S(_09335_),
    .X(_09339_));
 sky130_fd_sc_hd__buf_2 _15773_ (.A(_09339_),
    .X(_09340_));
 sky130_fd_sc_hd__clkbuf_4 _15774_ (.A(_09330_),
    .X(_09341_));
 sky130_fd_sc_hd__mux2_1 _15775_ (.A0(\core.cpuregs[23][2] ),
    .A1(_09340_),
    .S(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__buf_1 _15776_ (.A(_09342_),
    .X(_00278_));
 sky130_fd_sc_hd__buf_2 _15777_ (.A(_09334_),
    .X(_09343_));
 sky130_fd_sc_hd__nand2_1 _15778_ (.A(\core.reg_pc[3] ),
    .B(\core.reg_pc[2] ),
    .Y(_09344_));
 sky130_fd_sc_hd__inv_2 _15779_ (.A(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__nor2_1 _15780_ (.A(_09345_),
    .B(_09335_),
    .Y(_09346_));
 sky130_fd_sc_hd__or2_1 _15781_ (.A(\core.reg_pc[3] ),
    .B(\core.reg_pc[2] ),
    .X(_09347_));
 sky130_fd_sc_hd__a22o_1 _15782_ (.A1(_06641_),
    .A2(_09343_),
    .B1(_09346_),
    .B2(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__clkbuf_2 _15783_ (.A(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__mux2_1 _15784_ (.A0(\core.cpuregs[23][3] ),
    .A1(_09349_),
    .S(_09341_),
    .X(_09350_));
 sky130_fd_sc_hd__buf_1 _15785_ (.A(_09350_),
    .X(_00279_));
 sky130_fd_sc_hd__inv_2 _15786_ (.A(_09311_),
    .Y(_09351_));
 sky130_fd_sc_hd__clkbuf_2 _15787_ (.A(_09351_),
    .X(_09352_));
 sky130_fd_sc_hd__nand2_2 _15788_ (.A(_09345_),
    .B(\core.reg_pc[4] ),
    .Y(_09353_));
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(_09344_),
    .B(_07965_),
    .Y(_09354_));
 sky130_fd_sc_hd__and2_1 _15790_ (.A(_06669_),
    .B(_09312_),
    .X(_09355_));
 sky130_fd_sc_hd__a31o_2 _15791_ (.A1(_09352_),
    .A2(_09353_),
    .A3(_09354_),
    .B1(_09355_),
    .X(_09356_));
 sky130_fd_sc_hd__buf_2 _15792_ (.A(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__mux2_1 _15793_ (.A0(\core.cpuregs[23][4] ),
    .A1(_09357_),
    .S(_09341_),
    .X(_09358_));
 sky130_fd_sc_hd__buf_1 _15794_ (.A(_09358_),
    .X(_00280_));
 sky130_fd_sc_hd__nor2_2 _15795_ (.A(_08018_),
    .B(_09353_),
    .Y(_09359_));
 sky130_fd_sc_hd__nor2_1 _15796_ (.A(_09335_),
    .B(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(_09353_),
    .B(_08018_),
    .Y(_09361_));
 sky130_fd_sc_hd__a22o_1 _15798_ (.A1(_06695_),
    .A2(_09343_),
    .B1(_09360_),
    .B2(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__buf_2 _15799_ (.A(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(\core.cpuregs[23][5] ),
    .A1(_09363_),
    .S(_09341_),
    .X(_09364_));
 sky130_fd_sc_hd__clkbuf_1 _15801_ (.A(_09364_),
    .X(_00281_));
 sky130_fd_sc_hd__or2_1 _15802_ (.A(_05122_),
    .B(_09359_),
    .X(_09365_));
 sky130_fd_sc_hd__nand2_2 _15803_ (.A(_09359_),
    .B(_05122_),
    .Y(_09366_));
 sky130_fd_sc_hd__and2_1 _15804_ (.A(_06715_),
    .B(_09312_),
    .X(_09367_));
 sky130_fd_sc_hd__a31o_1 _15805_ (.A1(_09365_),
    .A2(_09352_),
    .A3(_09366_),
    .B1(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__buf_2 _15806_ (.A(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__mux2_1 _15807_ (.A0(\core.cpuregs[23][6] ),
    .A1(_09369_),
    .S(_09341_),
    .X(_09370_));
 sky130_fd_sc_hd__clkbuf_2 _15808_ (.A(_09370_),
    .X(_00282_));
 sky130_fd_sc_hd__or2_1 _15809_ (.A(_08112_),
    .B(_09366_),
    .X(_09371_));
 sky130_fd_sc_hd__nand2_2 _15810_ (.A(_09366_),
    .B(_08112_),
    .Y(_09372_));
 sky130_fd_sc_hd__and2_1 _15811_ (.A(_06734_),
    .B(_09312_),
    .X(_09373_));
 sky130_fd_sc_hd__a31o_1 _15812_ (.A1(_09371_),
    .A2(_09352_),
    .A3(_09372_),
    .B1(_09373_),
    .X(_09374_));
 sky130_fd_sc_hd__clkbuf_2 _15813_ (.A(_09374_),
    .X(_09375_));
 sky130_fd_sc_hd__mux2_1 _15814_ (.A0(\core.cpuregs[23][7] ),
    .A1(_09375_),
    .S(_09341_),
    .X(_09376_));
 sky130_fd_sc_hd__buf_1 _15815_ (.A(_09376_),
    .X(_00283_));
 sky130_fd_sc_hd__or2_1 _15816_ (.A(_08156_),
    .B(_09371_),
    .X(_09377_));
 sky130_fd_sc_hd__nand2_1 _15817_ (.A(_09371_),
    .B(_08156_),
    .Y(_09378_));
 sky130_fd_sc_hd__and2_1 _15818_ (.A(_06757_),
    .B(_09334_),
    .X(_09379_));
 sky130_fd_sc_hd__a31o_1 _15819_ (.A1(_09377_),
    .A2(_09351_),
    .A3(_09378_),
    .B1(_09379_),
    .X(_09380_));
 sky130_fd_sc_hd__clkbuf_2 _15820_ (.A(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(\core.cpuregs[23][8] ),
    .A1(_09381_),
    .S(_09330_),
    .X(_09382_));
 sky130_fd_sc_hd__clkbuf_1 _15822_ (.A(_09382_),
    .X(_00284_));
 sky130_fd_sc_hd__nand2_1 _15823_ (.A(_09377_),
    .B(_08203_),
    .Y(_09383_));
 sky130_fd_sc_hd__and4_1 _15824_ (.A(\core.reg_pc[9] ),
    .B(\core.reg_pc[8] ),
    .C(\core.reg_pc[7] ),
    .D(_05122_),
    .X(_09384_));
 sky130_fd_sc_hd__nand2_1 _15825_ (.A(_09384_),
    .B(_09359_),
    .Y(_09385_));
 sky130_fd_sc_hd__and2_1 _15826_ (.A(_06778_),
    .B(_09334_),
    .X(_09386_));
 sky130_fd_sc_hd__a31o_4 _15827_ (.A1(_09383_),
    .A2(_09351_),
    .A3(_09385_),
    .B1(_09386_),
    .X(_09387_));
 sky130_fd_sc_hd__clkbuf_4 _15828_ (.A(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(\core.cpuregs[23][9] ),
    .A1(_09388_),
    .S(_09330_),
    .X(_09389_));
 sky130_fd_sc_hd__buf_1 _15830_ (.A(_09389_),
    .X(_00285_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(_08263_),
    .B(_09385_),
    .Y(_09390_));
 sky130_fd_sc_hd__inv_2 _15832_ (.A(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand2_1 _15833_ (.A(_09385_),
    .B(_08263_),
    .Y(_09392_));
 sky130_fd_sc_hd__and2_1 _15834_ (.A(_06807_),
    .B(_09334_),
    .X(_09393_));
 sky130_fd_sc_hd__a31o_1 _15835_ (.A1(_09391_),
    .A2(_09351_),
    .A3(_09392_),
    .B1(_09393_),
    .X(_09394_));
 sky130_fd_sc_hd__buf_1 _15836_ (.A(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__mux2_1 _15837_ (.A0(\core.cpuregs[23][10] ),
    .A1(_09395_),
    .S(_09330_),
    .X(_09396_));
 sky130_fd_sc_hd__buf_1 _15838_ (.A(_09396_),
    .X(_00286_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_08348_),
    .B(_09391_),
    .Y(_09397_));
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(_09391_),
    .B(_08348_),
    .Y(_09398_));
 sky130_fd_sc_hd__or3b_1 _15841_ (.A(_09311_),
    .B(_09397_),
    .C_N(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__a21bo_1 _15842_ (.A1(_06829_),
    .A2(_09313_),
    .B1_N(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__buf_1 _15843_ (.A(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__inv_2 _15844_ (.A(_09329_),
    .Y(_09402_));
 sky130_fd_sc_hd__clkbuf_2 _15845_ (.A(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__mux2_1 _15846_ (.A0(_09401_),
    .A1(\core.cpuregs[23][11] ),
    .S(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__clkbuf_1 _15847_ (.A(_09404_),
    .X(_00287_));
 sky130_fd_sc_hd__o21a_1 _15848_ (.A1(\core.reg_pc[12] ),
    .A2(_09397_),
    .B1(_09351_),
    .X(_09405_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_09397_),
    .B(\core.reg_pc[12] ),
    .Y(_09406_));
 sky130_fd_sc_hd__a22o_1 _15850_ (.A1(_06854_),
    .A2(_09343_),
    .B1(_09405_),
    .B2(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__clkbuf_2 _15851_ (.A(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__mux2_2 _15852_ (.A0(\core.cpuregs[23][12] ),
    .A1(_09408_),
    .S(_09330_),
    .X(_09409_));
 sky130_fd_sc_hd__clkbuf_1 _15853_ (.A(_09409_),
    .X(_00288_));
 sky130_fd_sc_hd__and2_1 _15854_ (.A(_09406_),
    .B(_08447_),
    .X(_09410_));
 sky130_fd_sc_hd__nor2_4 _15855_ (.A(_08447_),
    .B(_09406_),
    .Y(_09411_));
 sky130_fd_sc_hd__or2_1 _15856_ (.A(_09311_),
    .B(_09411_),
    .X(_09412_));
 sky130_fd_sc_hd__a2bb2o_1 _15857_ (.A1_N(_09410_),
    .A2_N(_09412_),
    .B1(_06878_),
    .B2(_09343_),
    .X(_09413_));
 sky130_fd_sc_hd__clkbuf_2 _15858_ (.A(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__mux2_4 _15859_ (.A0(_09414_),
    .A1(\core.cpuregs[23][13] ),
    .S(_09403_),
    .X(_09415_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15860_ (.A(_09415_),
    .X(_00289_));
 sky130_fd_sc_hd__a21oi_1 _15861_ (.A1(_09411_),
    .A2(_07355_),
    .B1(_09335_),
    .Y(_09416_));
 sky130_fd_sc_hd__or2_1 _15862_ (.A(_07355_),
    .B(_09411_),
    .X(_09417_));
 sky130_fd_sc_hd__a22o_1 _15863_ (.A1(_06907_),
    .A2(_09343_),
    .B1(_09416_),
    .B2(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__buf_1 _15864_ (.A(_09418_),
    .X(_09419_));
 sky130_fd_sc_hd__mux2_1 _15865_ (.A0(_09419_),
    .A1(\core.cpuregs[23][14] ),
    .S(_09402_),
    .X(_09420_));
 sky130_fd_sc_hd__clkbuf_1 _15866_ (.A(_09420_),
    .X(_00290_));
 sky130_fd_sc_hd__a21oi_1 _15867_ (.A1(_09411_),
    .A2(_07355_),
    .B1(_05275_),
    .Y(_09421_));
 sky130_fd_sc_hd__a31o_1 _15868_ (.A1(_09411_),
    .A2(_05275_),
    .A3(_07355_),
    .B1(_09334_),
    .X(_09422_));
 sky130_fd_sc_hd__a2bb2o_1 _15869_ (.A1_N(_09421_),
    .A2_N(_09422_),
    .B1(_06930_),
    .B2(_09343_),
    .X(_09423_));
 sky130_fd_sc_hd__buf_1 _15870_ (.A(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__mux2_4 _15871_ (.A0(_09424_),
    .A1(\core.cpuregs[23][15] ),
    .S(_09402_),
    .X(_09425_));
 sky130_fd_sc_hd__clkbuf_1 _15872_ (.A(_09425_),
    .X(_00291_));
 sky130_fd_sc_hd__nand2_2 _15873_ (.A(_05275_),
    .B(\core.reg_pc[14] ),
    .Y(_09426_));
 sky130_fd_sc_hd__or4_1 _15874_ (.A(_08447_),
    .B(_08396_),
    .C(_08348_),
    .D(_08263_),
    .X(_09427_));
 sky130_fd_sc_hd__nor3_1 _15875_ (.A(_09385_),
    .B(_09426_),
    .C(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__xor2_1 _15876_ (.A(\core.reg_pc[16] ),
    .B(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__mux2_4 _15877_ (.A0(_09429_),
    .A1(_06962_),
    .S(_09312_),
    .X(_09430_));
 sky130_fd_sc_hd__buf_1 _15878_ (.A(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__mux2_1 _15879_ (.A0(_09431_),
    .A1(\core.cpuregs[23][16] ),
    .S(_09402_),
    .X(_09432_));
 sky130_fd_sc_hd__clkbuf_1 _15880_ (.A(_09432_),
    .X(_00292_));
 sky130_fd_sc_hd__nand2_1 _15881_ (.A(_09428_),
    .B(\core.reg_pc[16] ),
    .Y(_09433_));
 sky130_fd_sc_hd__xor2_1 _15882_ (.A(_08657_),
    .B(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__mux2_1 _15883_ (.A0(_09434_),
    .A1(_06984_),
    .S(_09312_),
    .X(_09435_));
 sky130_fd_sc_hd__buf_2 _15884_ (.A(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__mux2_1 _15885_ (.A0(_09436_),
    .A1(\core.cpuregs[23][17] ),
    .S(_09402_),
    .X(_09437_));
 sky130_fd_sc_hd__clkbuf_1 _15886_ (.A(_09437_),
    .X(_00293_));
 sky130_fd_sc_hd__or4_1 _15887_ (.A(_08657_),
    .B(_08610_),
    .C(_09426_),
    .D(_09427_),
    .X(_09438_));
 sky130_fd_sc_hd__nor2_1 _15888_ (.A(_09385_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__xor2_1 _15889_ (.A(_05339_),
    .B(_09439_),
    .X(_09440_));
 sky130_fd_sc_hd__mux2_1 _15890_ (.A0(_09440_),
    .A1(_07017_),
    .S(_09313_),
    .X(_09441_));
 sky130_fd_sc_hd__clkbuf_2 _15891_ (.A(_09441_),
    .X(_09442_));
 sky130_fd_sc_hd__nand2_1 _15892_ (.A(_09403_),
    .B(\core.cpuregs[23][18] ),
    .Y(_09443_));
 sky130_fd_sc_hd__a21bo_1 _15893_ (.A1(_09442_),
    .A2(_09331_),
    .B1_N(_09443_),
    .X(_00294_));
 sky130_fd_sc_hd__nand2_1 _15894_ (.A(_09439_),
    .B(_05339_),
    .Y(_09444_));
 sky130_fd_sc_hd__xor2_1 _15895_ (.A(_08759_),
    .B(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__clkbuf_4 _15896_ (.A(_09335_),
    .X(_09446_));
 sky130_fd_sc_hd__mux2_4 _15897_ (.A0(_09445_),
    .A1(_07041_),
    .S(_09446_),
    .X(_09447_));
 sky130_fd_sc_hd__buf_4 _15898_ (.A(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__clkbuf_2 _15899_ (.A(_09331_),
    .X(_09449_));
 sky130_fd_sc_hd__nand2_2 _15900_ (.A(_09448_),
    .B(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__clkbuf_4 _15901_ (.A(_09403_),
    .X(_09451_));
 sky130_fd_sc_hd__nand2_1 _15902_ (.A(_09451_),
    .B(\core.cpuregs[23][19] ),
    .Y(_09452_));
 sky130_fd_sc_hd__nand2_2 _15903_ (.A(_09450_),
    .B(_09452_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_2 _15904_ (.A(\core.reg_pc[19] ),
    .B(\core.reg_pc[18] ),
    .Y(_09453_));
 sky130_fd_sc_hd__inv_2 _15905_ (.A(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_09439_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__xor2_1 _15907_ (.A(_08806_),
    .B(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__mux2_4 _15908_ (.A0(_09456_),
    .A1(_07067_),
    .S(_09446_),
    .X(_09457_));
 sky130_fd_sc_hd__clkbuf_2 _15909_ (.A(_09457_),
    .X(_09458_));
 sky130_fd_sc_hd__nand2_1 _15910_ (.A(_09458_),
    .B(_09449_),
    .Y(_09459_));
 sky130_fd_sc_hd__nand2_1 _15911_ (.A(_09451_),
    .B(\core.cpuregs[23][20] ),
    .Y(_09460_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_09459_),
    .B(_09460_),
    .Y(_00296_));
 sky130_fd_sc_hd__buf_4 _15913_ (.A(_09313_),
    .X(_09461_));
 sky130_fd_sc_hd__or2_1 _15914_ (.A(_08806_),
    .B(_09455_),
    .X(_09462_));
 sky130_fd_sc_hd__xor2_2 _15915_ (.A(\core.reg_pc[21] ),
    .B(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__clkbuf_4 _15916_ (.A(_09313_),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_1 _15917_ (.A(_07090_),
    .B(_09464_),
    .Y(_09465_));
 sky130_fd_sc_hd__o21ai_4 _15918_ (.A1(_09461_),
    .A2(_09463_),
    .B1(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__buf_6 _15919_ (.A(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__nand2_1 _15920_ (.A(_09467_),
    .B(_09449_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_1 _15921_ (.A(_09451_),
    .B(\core.cpuregs[23][21] ),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_1 _15922_ (.A(_09468_),
    .B(_09469_),
    .Y(_00297_));
 sky130_fd_sc_hd__and3_1 _15923_ (.A(_09454_),
    .B(\core.reg_pc[21] ),
    .C(\core.reg_pc[20] ),
    .X(_09470_));
 sky130_fd_sc_hd__nand2_2 _15924_ (.A(_09439_),
    .B(_09470_),
    .Y(_09471_));
 sky130_fd_sc_hd__xor2_1 _15925_ (.A(_08914_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__mux2_1 _15926_ (.A0(_09472_),
    .A1(_07119_),
    .S(_09313_),
    .X(_09473_));
 sky130_fd_sc_hd__clkbuf_2 _15927_ (.A(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(_09474_),
    .B(_09449_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand2_1 _15929_ (.A(_09451_),
    .B(\core.cpuregs[23][22] ),
    .Y(_09476_));
 sky130_fd_sc_hd__nand2_1 _15930_ (.A(_09475_),
    .B(_09476_),
    .Y(_00298_));
 sky130_fd_sc_hd__or2_1 _15931_ (.A(_08914_),
    .B(_09471_),
    .X(_09477_));
 sky130_fd_sc_hd__xor2_2 _15932_ (.A(\core.reg_pc[23] ),
    .B(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(_07138_),
    .B(_09464_),
    .Y(_09479_));
 sky130_fd_sc_hd__o21ai_4 _15934_ (.A1(_09461_),
    .A2(_09478_),
    .B1(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__buf_6 _15935_ (.A(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__nand2_1 _15936_ (.A(_09481_),
    .B(_09449_),
    .Y(_09482_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(_09451_),
    .B(\core.cpuregs[23][23] ),
    .Y(_09483_));
 sky130_fd_sc_hd__nand2_1 _15938_ (.A(_09482_),
    .B(_09483_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _15939_ (.A(\core.reg_pc[23] ),
    .B(\core.reg_pc[22] ),
    .Y(_09484_));
 sky130_fd_sc_hd__or2_1 _15940_ (.A(_09484_),
    .B(_09471_),
    .X(_09485_));
 sky130_fd_sc_hd__xor2_2 _15941_ (.A(\core.reg_pc[24] ),
    .B(_09485_),
    .X(_09486_));
 sky130_fd_sc_hd__nand2_1 _15942_ (.A(_07162_),
    .B(_09464_),
    .Y(_09487_));
 sky130_fd_sc_hd__o21ai_4 _15943_ (.A1(_09461_),
    .A2(_09486_),
    .B1(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__buf_6 _15944_ (.A(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__nand2_4 _15945_ (.A(_09489_),
    .B(_09449_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(_09451_),
    .B(\core.cpuregs[23][24] ),
    .Y(_09491_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(_09490_),
    .B(_09491_),
    .Y(_00300_));
 sky130_fd_sc_hd__o21ai_1 _15948_ (.A1(_09005_),
    .A2(_09485_),
    .B1(\core.reg_pc[25] ),
    .Y(_09492_));
 sky130_fd_sc_hd__nor2_1 _15949_ (.A(_09005_),
    .B(_09485_),
    .Y(_09493_));
 sky130_fd_sc_hd__nand2_1 _15950_ (.A(_09493_),
    .B(_09052_),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_1 _15951_ (.A(_09492_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__nand2_1 _15952_ (.A(_09495_),
    .B(_09352_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(_07185_),
    .B(_09461_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand2_1 _15954_ (.A(_09496_),
    .B(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__buf_2 _15955_ (.A(_09498_),
    .X(_09499_));
 sky130_fd_sc_hd__clkbuf_4 _15956_ (.A(_09331_),
    .X(_09500_));
 sky130_fd_sc_hd__nand2_4 _15957_ (.A(_09499_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15958_ (.A(_09403_),
    .X(_09502_));
 sky130_fd_sc_hd__nand2_1 _15959_ (.A(_09502_),
    .B(\core.cpuregs[23][25] ),
    .Y(_09503_));
 sky130_fd_sc_hd__nand2_1 _15960_ (.A(_09501_),
    .B(_09503_),
    .Y(_00301_));
 sky130_fd_sc_hd__and4b_1 _15961_ (.A_N(_09484_),
    .B(_09470_),
    .C(\core.reg_pc[25] ),
    .D(\core.reg_pc[24] ),
    .X(_09504_));
 sky130_fd_sc_hd__and2_1 _15962_ (.A(_09439_),
    .B(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__buf_6 _15963_ (.A(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__xor2_2 _15964_ (.A(_05464_),
    .B(_09506_),
    .X(_09507_));
 sky130_fd_sc_hd__mux2_1 _15965_ (.A0(_09507_),
    .A1(_07216_),
    .S(_09446_),
    .X(_09508_));
 sky130_fd_sc_hd__clkbuf_4 _15966_ (.A(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__nand2_1 _15967_ (.A(_09509_),
    .B(_09500_),
    .Y(_09510_));
 sky130_fd_sc_hd__nand2_2 _15968_ (.A(_09502_),
    .B(\core.cpuregs[23][26] ),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_1 _15969_ (.A(_09510_),
    .B(_09511_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _15970_ (.A(_09506_),
    .B(_05464_),
    .Y(_09512_));
 sky130_fd_sc_hd__xor2_2 _15971_ (.A(\core.reg_pc[27] ),
    .B(_09512_),
    .X(_09513_));
 sky130_fd_sc_hd__nand2_1 _15972_ (.A(_07234_),
    .B(_09464_),
    .Y(_09514_));
 sky130_fd_sc_hd__o21ai_4 _15973_ (.A1(_09446_),
    .A2(_09513_),
    .B1(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__buf_6 _15974_ (.A(_09515_),
    .X(_09516_));
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(_09516_),
    .B(_09500_),
    .Y(_09517_));
 sky130_fd_sc_hd__nand2_1 _15976_ (.A(_09502_),
    .B(\core.cpuregs[23][27] ),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_1 _15977_ (.A(_09517_),
    .B(_09518_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _15978_ (.A(\core.reg_pc[27] ),
    .B(\core.reg_pc[26] ),
    .Y(_09519_));
 sky130_fd_sc_hd__inv_2 _15979_ (.A(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_2 _15980_ (.A(_09506_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__xor2_2 _15981_ (.A(_05492_),
    .B(_09521_),
    .X(_09522_));
 sky130_fd_sc_hd__nand2_1 _15982_ (.A(_07256_),
    .B(_09464_),
    .Y(_09523_));
 sky130_fd_sc_hd__o21ai_4 _15983_ (.A1(_09446_),
    .A2(_09522_),
    .B1(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__buf_6 _15984_ (.A(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__nand2_1 _15985_ (.A(_09525_),
    .B(_09500_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand2_1 _15986_ (.A(_09502_),
    .B(\core.cpuregs[23][28] ),
    .Y(_09527_));
 sky130_fd_sc_hd__nand2_1 _15987_ (.A(_09526_),
    .B(_09527_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand3b_1 _15988_ (.A_N(_09521_),
    .B(_09237_),
    .C(_05492_),
    .Y(_09528_));
 sky130_fd_sc_hd__o21ai_1 _15989_ (.A1(_09193_),
    .A2(_09521_),
    .B1(\core.reg_pc[29] ),
    .Y(_09529_));
 sky130_fd_sc_hd__nand2_1 _15990_ (.A(_09528_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__nand2_1 _15991_ (.A(_09530_),
    .B(_09352_),
    .Y(_09531_));
 sky130_fd_sc_hd__nand2_1 _15992_ (.A(_07282_),
    .B(_09461_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__buf_4 _15994_ (.A(_09533_),
    .X(_09534_));
 sky130_fd_sc_hd__nand2_1 _15995_ (.A(_09534_),
    .B(_09500_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_1 _15996_ (.A(_09502_),
    .B(\core.cpuregs[23][29] ),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_1 _15997_ (.A(_09535_),
    .B(_09536_),
    .Y(_00305_));
 sky130_fd_sc_hd__and3_1 _15998_ (.A(_09520_),
    .B(\core.reg_pc[29] ),
    .C(\core.reg_pc[28] ),
    .X(_09537_));
 sky130_fd_sc_hd__nand2_2 _15999_ (.A(_09506_),
    .B(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__xor2_2 _16000_ (.A(\core.reg_pc[30] ),
    .B(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__nand2_1 _16001_ (.A(_07308_),
    .B(_09464_),
    .Y(_09540_));
 sky130_fd_sc_hd__o21ai_4 _16002_ (.A1(_09446_),
    .A2(_09539_),
    .B1(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__buf_6 _16003_ (.A(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__nand2_1 _16004_ (.A(_09542_),
    .B(_09500_),
    .Y(_09543_));
 sky130_fd_sc_hd__nand2_1 _16005_ (.A(_09502_),
    .B(\core.cpuregs[23][30] ),
    .Y(_09544_));
 sky130_fd_sc_hd__nand2_1 _16006_ (.A(_09543_),
    .B(_09544_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand3b_1 _16007_ (.A_N(_09538_),
    .B(_06303_),
    .C(\core.reg_pc[30] ),
    .Y(_09545_));
 sky130_fd_sc_hd__o21ai_1 _16008_ (.A1(_05518_),
    .A2(_09538_),
    .B1(\core.reg_pc[31] ),
    .Y(_09546_));
 sky130_fd_sc_hd__nand2_1 _16009_ (.A(_09545_),
    .B(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__nand2_1 _16010_ (.A(_09547_),
    .B(_09352_),
    .Y(_09548_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(_07334_),
    .B(_09461_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_1 _16012_ (.A(_09548_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__clkbuf_2 _16013_ (.A(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__nand2_1 _16014_ (.A(_09551_),
    .B(_09331_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand2_1 _16015_ (.A(_09403_),
    .B(\core.cpuregs[23][31] ),
    .Y(_09553_));
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(_09552_),
    .B(_09553_),
    .Y(_00307_));
 sky130_fd_sc_hd__buf_1 _16017_ (.A(_09323_),
    .X(_09554_));
 sky130_fd_sc_hd__inv_2 _16018_ (.A(\core.latched_rd[1] ),
    .Y(_09555_));
 sky130_fd_sc_hd__nor2_1 _16019_ (.A(\core.latched_rd[0] ),
    .B(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__and3_1 _16020_ (.A(\core.latched_rd[4] ),
    .B(\core.latched_rd[3] ),
    .C(\core.latched_rd[2] ),
    .X(_09557_));
 sky130_fd_sc_hd__and3_2 _16021_ (.A(_09554_),
    .B(_09556_),
    .C(_09557_),
    .X(_09558_));
 sky130_fd_sc_hd__clkbuf_2 _16022_ (.A(_09558_),
    .X(_09559_));
 sky130_fd_sc_hd__clkbuf_2 _16023_ (.A(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__mux2_1 _16024_ (.A0(\core.cpuregs[30][0] ),
    .A1(_09315_),
    .S(_09560_),
    .X(_09561_));
 sky130_fd_sc_hd__buf_1 _16025_ (.A(_09561_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_2 _16026_ (.A0(\core.cpuregs[30][1] ),
    .A1(_09337_),
    .S(_09560_),
    .X(_09562_));
 sky130_fd_sc_hd__clkbuf_1 _16027_ (.A(_09562_),
    .X(_00309_));
 sky130_fd_sc_hd__clkbuf_4 _16028_ (.A(_09559_),
    .X(_09563_));
 sky130_fd_sc_hd__mux2_1 _16029_ (.A0(\core.cpuregs[30][2] ),
    .A1(_09340_),
    .S(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__clkbuf_1 _16030_ (.A(_09564_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _16031_ (.A0(\core.cpuregs[30][3] ),
    .A1(_09349_),
    .S(_09563_),
    .X(_09565_));
 sky130_fd_sc_hd__buf_1 _16032_ (.A(_09565_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _16033_ (.A0(\core.cpuregs[30][4] ),
    .A1(_09357_),
    .S(_09563_),
    .X(_09566_));
 sky130_fd_sc_hd__buf_1 _16034_ (.A(_09566_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _16035_ (.A0(\core.cpuregs[30][5] ),
    .A1(_09363_),
    .S(_09563_),
    .X(_09567_));
 sky130_fd_sc_hd__clkbuf_1 _16036_ (.A(_09567_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _16037_ (.A0(\core.cpuregs[30][6] ),
    .A1(_09369_),
    .S(_09563_),
    .X(_09568_));
 sky130_fd_sc_hd__clkbuf_1 _16038_ (.A(_09568_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _16039_ (.A0(\core.cpuregs[30][7] ),
    .A1(_09375_),
    .S(_09563_),
    .X(_09569_));
 sky130_fd_sc_hd__clkbuf_1 _16040_ (.A(_09569_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _16041_ (.A0(\core.cpuregs[30][8] ),
    .A1(_09381_),
    .S(_09559_),
    .X(_09570_));
 sky130_fd_sc_hd__clkbuf_1 _16042_ (.A(_09570_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _16043_ (.A0(\core.cpuregs[30][9] ),
    .A1(_09388_),
    .S(_09559_),
    .X(_09571_));
 sky130_fd_sc_hd__clkbuf_1 _16044_ (.A(_09571_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _16045_ (.A0(\core.cpuregs[30][10] ),
    .A1(_09395_),
    .S(_09559_),
    .X(_09572_));
 sky130_fd_sc_hd__buf_1 _16046_ (.A(_09572_),
    .X(_00318_));
 sky130_fd_sc_hd__inv_2 _16047_ (.A(_09558_),
    .Y(_09573_));
 sky130_fd_sc_hd__clkbuf_2 _16048_ (.A(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__mux2_1 _16049_ (.A0(_09401_),
    .A1(\core.cpuregs[30][11] ),
    .S(_09574_),
    .X(_09575_));
 sky130_fd_sc_hd__clkbuf_1 _16050_ (.A(_09575_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_8 _16051_ (.A0(\core.cpuregs[30][12] ),
    .A1(_09408_),
    .S(_09559_),
    .X(_09576_));
 sky130_fd_sc_hd__clkbuf_1 _16052_ (.A(_09576_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _16053_ (.A0(_09414_),
    .A1(\core.cpuregs[30][13] ),
    .S(_09574_),
    .X(_09577_));
 sky130_fd_sc_hd__buf_1 _16054_ (.A(_09577_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_4 _16055_ (.A0(_09419_),
    .A1(\core.cpuregs[30][14] ),
    .S(_09573_),
    .X(_09578_));
 sky130_fd_sc_hd__clkbuf_1 _16056_ (.A(_09578_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _16057_ (.A0(_09424_),
    .A1(\core.cpuregs[30][15] ),
    .S(_09573_),
    .X(_09579_));
 sky130_fd_sc_hd__clkbuf_1 _16058_ (.A(_09579_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _16059_ (.A0(_09431_),
    .A1(\core.cpuregs[30][16] ),
    .S(_09573_),
    .X(_09580_));
 sky130_fd_sc_hd__clkbuf_1 _16060_ (.A(_09580_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _16061_ (.A0(_09436_),
    .A1(\core.cpuregs[30][17] ),
    .S(_09573_),
    .X(_09581_));
 sky130_fd_sc_hd__clkbuf_1 _16062_ (.A(_09581_),
    .X(_00325_));
 sky130_fd_sc_hd__nand2_1 _16063_ (.A(_09574_),
    .B(\core.cpuregs[30][18] ),
    .Y(_09582_));
 sky130_fd_sc_hd__a21bo_1 _16064_ (.A1(_09442_),
    .A2(_09560_),
    .B1_N(_09582_),
    .X(_00326_));
 sky130_fd_sc_hd__clkbuf_2 _16065_ (.A(_09560_),
    .X(_09583_));
 sky130_fd_sc_hd__nand2_1 _16066_ (.A(_09448_),
    .B(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__buf_4 _16067_ (.A(_09574_),
    .X(_09585_));
 sky130_fd_sc_hd__nand2_2 _16068_ (.A(_09585_),
    .B(\core.cpuregs[30][19] ),
    .Y(_09586_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(_09584_),
    .B(_09586_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_4 _16070_ (.A(_09458_),
    .B(_09583_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand2_4 _16071_ (.A(_09585_),
    .B(\core.cpuregs[30][20] ),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_1 _16072_ (.A(_09587_),
    .B(_09588_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(_09467_),
    .B(_09583_),
    .Y(_09589_));
 sky130_fd_sc_hd__nand2_1 _16074_ (.A(_09585_),
    .B(\core.cpuregs[30][21] ),
    .Y(_09590_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(_09589_),
    .B(_09590_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_2 _16076_ (.A(_09474_),
    .B(_09583_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand2_4 _16077_ (.A(_09585_),
    .B(\core.cpuregs[30][22] ),
    .Y(_09592_));
 sky130_fd_sc_hd__nand2_1 _16078_ (.A(_09591_),
    .B(_09592_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _16079_ (.A(_09481_),
    .B(_09583_),
    .Y(_09593_));
 sky130_fd_sc_hd__nand2_1 _16080_ (.A(_09585_),
    .B(\core.cpuregs[30][23] ),
    .Y(_09594_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(_09593_),
    .B(_09594_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _16082_ (.A(_09489_),
    .B(_09583_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(_09585_),
    .B(\core.cpuregs[30][24] ),
    .Y(_09596_));
 sky130_fd_sc_hd__nand2_1 _16084_ (.A(_09595_),
    .B(_09596_),
    .Y(_00332_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16085_ (.A(_09560_),
    .X(_09597_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_09499_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__clkbuf_2 _16087_ (.A(_09574_),
    .X(_09599_));
 sky130_fd_sc_hd__nand2_2 _16088_ (.A(_09599_),
    .B(\core.cpuregs[30][25] ),
    .Y(_09600_));
 sky130_fd_sc_hd__nand2_2 _16089_ (.A(_09598_),
    .B(_09600_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _16090_ (.A(_09509_),
    .B(_09597_),
    .Y(_09601_));
 sky130_fd_sc_hd__nand2_1 _16091_ (.A(_09599_),
    .B(\core.cpuregs[30][26] ),
    .Y(_09602_));
 sky130_fd_sc_hd__nand2_1 _16092_ (.A(_09601_),
    .B(_09602_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _16093_ (.A(_09516_),
    .B(_09597_),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_1 _16094_ (.A(_09599_),
    .B(\core.cpuregs[30][27] ),
    .Y(_09604_));
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(_09603_),
    .B(_09604_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _16096_ (.A(_09525_),
    .B(_09597_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(_09599_),
    .B(\core.cpuregs[30][28] ),
    .Y(_09606_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(_09605_),
    .B(_09606_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(_09534_),
    .B(_09597_),
    .Y(_09607_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(_09599_),
    .B(net117),
    .Y(_09608_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(_09607_),
    .B(_09608_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _16102_ (.A(_09542_),
    .B(_09597_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_2 _16103_ (.A(_09599_),
    .B(\core.cpuregs[30][30] ),
    .Y(_09610_));
 sky130_fd_sc_hd__nand2_1 _16104_ (.A(_09609_),
    .B(_09610_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(_09551_),
    .B(_09560_),
    .Y(_09611_));
 sky130_fd_sc_hd__nand2_2 _16106_ (.A(_09574_),
    .B(\core.cpuregs[30][31] ),
    .Y(_09612_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(_09611_),
    .B(_09612_),
    .Y(_00339_));
 sky130_fd_sc_hd__clkbuf_2 _16108_ (.A(_04520_),
    .X(_09613_));
 sky130_fd_sc_hd__mux2_1 _16109_ (.A0(\core.cpuregs[0][0] ),
    .A1(\core.cpuregs[1][0] ),
    .S(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__clkbuf_2 _16110_ (.A(_04524_),
    .X(_09615_));
 sky130_fd_sc_hd__mux2_1 _16111_ (.A0(\core.cpuregs[2][0] ),
    .A1(\core.cpuregs[3][0] ),
    .S(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__clkbuf_2 _16112_ (.A(_04640_),
    .X(_09617_));
 sky130_fd_sc_hd__mux2_1 _16113_ (.A0(_09614_),
    .A1(_09616_),
    .S(_09617_),
    .X(_09618_));
 sky130_fd_sc_hd__mux2_1 _16114_ (.A0(\core.cpuregs[6][0] ),
    .A1(\core.cpuregs[7][0] ),
    .S(_09613_),
    .X(_09619_));
 sky130_fd_sc_hd__clkbuf_2 _16115_ (.A(_04524_),
    .X(_09620_));
 sky130_fd_sc_hd__mux2_1 _16116_ (.A0(\core.cpuregs[4][0] ),
    .A1(\core.cpuregs[5][0] ),
    .S(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__clkbuf_2 _16117_ (.A(_04536_),
    .X(_09622_));
 sky130_fd_sc_hd__mux2_1 _16118_ (.A0(_09619_),
    .A1(_09621_),
    .S(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__clkbuf_2 _16119_ (.A(_00002_),
    .X(_09624_));
 sky130_fd_sc_hd__mux2_1 _16120_ (.A0(_09618_),
    .A1(_09623_),
    .S(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__mux2_1 _16121_ (.A0(\core.cpuregs[12][0] ),
    .A1(\core.cpuregs[13][0] ),
    .S(_09613_),
    .X(_09626_));
 sky130_fd_sc_hd__mux2_1 _16122_ (.A0(\core.cpuregs[14][0] ),
    .A1(\core.cpuregs[15][0] ),
    .S(_09620_),
    .X(_09627_));
 sky130_fd_sc_hd__mux2_1 _16123_ (.A0(_09626_),
    .A1(_09627_),
    .S(_09617_),
    .X(_09628_));
 sky130_fd_sc_hd__mux2_1 _16124_ (.A0(\core.cpuregs[8][0] ),
    .A1(\core.cpuregs[9][0] ),
    .S(_09615_),
    .X(_09629_));
 sky130_fd_sc_hd__clkbuf_2 _16125_ (.A(_04524_),
    .X(_09630_));
 sky130_fd_sc_hd__mux2_1 _16126_ (.A0(\core.cpuregs[10][0] ),
    .A1(\core.cpuregs[11][0] ),
    .S(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__clkbuf_2 _16127_ (.A(_04528_),
    .X(_09632_));
 sky130_fd_sc_hd__mux2_1 _16128_ (.A0(_09629_),
    .A1(_09631_),
    .S(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__mux2_1 _16129_ (.A0(_09628_),
    .A1(_09633_),
    .S(_04550_),
    .X(_09634_));
 sky130_fd_sc_hd__mux2_1 _16130_ (.A0(_09625_),
    .A1(_09634_),
    .S(_04656_),
    .X(_09635_));
 sky130_fd_sc_hd__mux2_1 _16131_ (.A0(\core.cpuregs[16][0] ),
    .A1(\core.cpuregs[17][0] ),
    .S(_09615_),
    .X(_09636_));
 sky130_fd_sc_hd__mux2_1 _16132_ (.A0(\core.cpuregs[18][0] ),
    .A1(\core.cpuregs[19][0] ),
    .S(_09630_),
    .X(_09637_));
 sky130_fd_sc_hd__mux2_1 _16133_ (.A0(_09636_),
    .A1(_09637_),
    .S(_09632_),
    .X(_09638_));
 sky130_fd_sc_hd__mux2_1 _16134_ (.A0(\core.cpuregs[22][0] ),
    .A1(\core.cpuregs[23][0] ),
    .S(_09630_),
    .X(_09639_));
 sky130_fd_sc_hd__clkbuf_2 _16135_ (.A(_04524_),
    .X(_09640_));
 sky130_fd_sc_hd__mux2_1 _16136_ (.A0(\core.cpuregs[20][0] ),
    .A1(\core.cpuregs[21][0] ),
    .S(_09640_),
    .X(_09641_));
 sky130_fd_sc_hd__mux2_1 _16137_ (.A0(_09639_),
    .A1(_09641_),
    .S(_09622_),
    .X(_09642_));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(_09638_),
    .A1(_09642_),
    .S(_09624_),
    .X(_09643_));
 sky130_fd_sc_hd__mux2_1 _16139_ (.A0(\core.cpuregs[24][0] ),
    .A1(\core.cpuregs[25][0] ),
    .S(_09620_),
    .X(_09644_));
 sky130_fd_sc_hd__mux2_4 _16140_ (.A0(\core.cpuregs[26][0] ),
    .A1(\core.cpuregs[27][0] ),
    .S(_09640_),
    .X(_09645_));
 sky130_fd_sc_hd__mux2_1 _16141_ (.A0(_09644_),
    .A1(_09645_),
    .S(_09632_),
    .X(_09646_));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(\core.cpuregs[28][0] ),
    .A1(\core.cpuregs[29][0] ),
    .S(_09640_),
    .X(_09647_));
 sky130_fd_sc_hd__clkbuf_2 _16143_ (.A(_04520_),
    .X(_09648_));
 sky130_fd_sc_hd__mux2_1 _16144_ (.A0(\core.cpuregs[30][0] ),
    .A1(\core.cpuregs[31][0] ),
    .S(_09648_),
    .X(_09649_));
 sky130_fd_sc_hd__clkbuf_2 _16145_ (.A(_04528_),
    .X(_09650_));
 sky130_fd_sc_hd__mux2_1 _16146_ (.A0(_09647_),
    .A1(_09649_),
    .S(_09650_),
    .X(_09651_));
 sky130_fd_sc_hd__mux2_1 _16147_ (.A0(_09646_),
    .A1(_09651_),
    .S(_09624_),
    .X(_09652_));
 sky130_fd_sc_hd__mux2_1 _16148_ (.A0(_09643_),
    .A1(_09652_),
    .S(_04656_),
    .X(_09653_));
 sky130_fd_sc_hd__mux2_1 _16149_ (.A0(_09635_),
    .A1(_09653_),
    .S(_04573_),
    .X(_09654_));
 sky130_fd_sc_hd__nand2_1 _16150_ (.A(_09654_),
    .B(_04582_),
    .Y(_09655_));
 sky130_fd_sc_hd__or2_1 _16151_ (.A(_04485_),
    .B(_09655_),
    .X(_09656_));
 sky130_fd_sc_hd__a21oi_1 _16152_ (.A1(_04577_),
    .A2(_04485_),
    .B1(_05063_),
    .Y(_09657_));
 sky130_fd_sc_hd__o21ai_1 _16153_ (.A1(\core.reg_sh[0] ),
    .A2(_07660_),
    .B1(_05115_),
    .Y(_09658_));
 sky130_fd_sc_hd__a21bo_1 _16154_ (.A1(_09656_),
    .A2(_09657_),
    .B1_N(_09658_),
    .X(_09659_));
 sky130_fd_sc_hd__nand2_1 _16155_ (.A(_04627_),
    .B(\core.reg_sh[0] ),
    .Y(_09660_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_09659_),
    .B(_09660_),
    .Y(_00340_));
 sky130_fd_sc_hd__mux2_1 _16157_ (.A0(\core.cpuregs[0][1] ),
    .A1(\core.cpuregs[1][1] ),
    .S(_09613_),
    .X(_09661_));
 sky130_fd_sc_hd__mux2_1 _16158_ (.A0(\core.cpuregs[2][1] ),
    .A1(\core.cpuregs[3][1] ),
    .S(_09615_),
    .X(_09662_));
 sky130_fd_sc_hd__mux2_1 _16159_ (.A0(_09661_),
    .A1(_09662_),
    .S(_09617_),
    .X(_09663_));
 sky130_fd_sc_hd__mux2_1 _16160_ (.A0(\core.cpuregs[6][1] ),
    .A1(\core.cpuregs[7][1] ),
    .S(_09615_),
    .X(_09664_));
 sky130_fd_sc_hd__mux2_1 _16161_ (.A0(\core.cpuregs[4][1] ),
    .A1(\core.cpuregs[5][1] ),
    .S(_09620_),
    .X(_09665_));
 sky130_fd_sc_hd__mux2_1 _16162_ (.A0(_09664_),
    .A1(_09665_),
    .S(_09622_),
    .X(_09666_));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(_09663_),
    .A1(_09666_),
    .S(_09624_),
    .X(_09667_));
 sky130_fd_sc_hd__mux2_1 _16164_ (.A0(\core.cpuregs[12][1] ),
    .A1(\core.cpuregs[13][1] ),
    .S(_09613_),
    .X(_09668_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(\core.cpuregs[14][1] ),
    .A1(\core.cpuregs[15][1] ),
    .S(_09620_),
    .X(_09669_));
 sky130_fd_sc_hd__mux2_1 _16166_ (.A0(_09668_),
    .A1(_09669_),
    .S(_09632_),
    .X(_09670_));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(\core.cpuregs[8][1] ),
    .A1(\core.cpuregs[9][1] ),
    .S(_09620_),
    .X(_09671_));
 sky130_fd_sc_hd__mux2_1 _16168_ (.A0(\core.cpuregs[10][1] ),
    .A1(\core.cpuregs[11][1] ),
    .S(_09640_),
    .X(_09672_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(_09671_),
    .A1(_09672_),
    .S(_09632_),
    .X(_09673_));
 sky130_fd_sc_hd__mux2_1 _16170_ (.A0(_09670_),
    .A1(_09673_),
    .S(_04550_),
    .X(_09674_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(_09667_),
    .A1(_09674_),
    .S(_04656_),
    .X(_09675_));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(\core.cpuregs[16][1] ),
    .A1(\core.cpuregs[17][1] ),
    .S(_09615_),
    .X(_09676_));
 sky130_fd_sc_hd__mux2_1 _16173_ (.A0(\core.cpuregs[18][1] ),
    .A1(\core.cpuregs[19][1] ),
    .S(_09630_),
    .X(_09677_));
 sky130_fd_sc_hd__mux2_1 _16174_ (.A0(_09676_),
    .A1(_09677_),
    .S(_09632_),
    .X(_09678_));
 sky130_fd_sc_hd__mux2_4 _16175_ (.A0(\core.cpuregs[22][1] ),
    .A1(\core.cpuregs[23][1] ),
    .S(_09630_),
    .X(_09679_));
 sky130_fd_sc_hd__mux2_1 _16176_ (.A0(\core.cpuregs[20][1] ),
    .A1(\core.cpuregs[21][1] ),
    .S(_09648_),
    .X(_09680_));
 sky130_fd_sc_hd__mux2_4 _16177_ (.A0(_09679_),
    .A1(_09680_),
    .S(_04536_),
    .X(_09681_));
 sky130_fd_sc_hd__mux2_1 _16178_ (.A0(_09678_),
    .A1(_09681_),
    .S(_09624_),
    .X(_09682_));
 sky130_fd_sc_hd__mux2_1 _16179_ (.A0(\core.cpuregs[24][1] ),
    .A1(\core.cpuregs[25][1] ),
    .S(_09630_),
    .X(_09683_));
 sky130_fd_sc_hd__mux2_1 _16180_ (.A0(\core.cpuregs[26][1] ),
    .A1(\core.cpuregs[27][1] ),
    .S(_09640_),
    .X(_09684_));
 sky130_fd_sc_hd__mux2_8 _16181_ (.A0(_09683_),
    .A1(_09684_),
    .S(_09650_),
    .X(_09685_));
 sky130_fd_sc_hd__mux2_1 _16182_ (.A0(\core.cpuregs[28][1] ),
    .A1(\core.cpuregs[29][1] ),
    .S(_09640_),
    .X(_09686_));
 sky130_fd_sc_hd__mux2_4 _16183_ (.A0(\core.cpuregs[30][1] ),
    .A1(\core.cpuregs[31][1] ),
    .S(_09648_),
    .X(_09687_));
 sky130_fd_sc_hd__mux2_1 _16184_ (.A0(_09686_),
    .A1(_09687_),
    .S(_09650_),
    .X(_09688_));
 sky130_fd_sc_hd__mux2_1 _16185_ (.A0(_09685_),
    .A1(_09688_),
    .S(_09624_),
    .X(_09689_));
 sky130_fd_sc_hd__mux2_1 _16186_ (.A0(_09682_),
    .A1(_09689_),
    .S(_00003_),
    .X(_09690_));
 sky130_fd_sc_hd__mux2_1 _16187_ (.A0(_09675_),
    .A1(_09690_),
    .S(_04573_),
    .X(_09691_));
 sky130_fd_sc_hd__nand2_1 _16188_ (.A(_09691_),
    .B(_04582_),
    .Y(_09692_));
 sky130_fd_sc_hd__or2_1 _16189_ (.A(\core.is_slli_srli_srai ),
    .B(_09692_),
    .X(_09693_));
 sky130_fd_sc_hd__a21oi_1 _16190_ (.A1(_05942_),
    .A2(_04485_),
    .B1(_05115_),
    .Y(_09694_));
 sky130_fd_sc_hd__or2b_1 _16191_ (.A(\core.reg_sh[1] ),
    .B_N(\core.reg_sh[0] ),
    .X(_09695_));
 sky130_fd_sc_hd__or2b_1 _16192_ (.A(\core.reg_sh[0] ),
    .B_N(\core.reg_sh[1] ),
    .X(_09696_));
 sky130_fd_sc_hd__a31o_1 _16193_ (.A1(_04589_),
    .A2(_09695_),
    .A3(_09696_),
    .B1(_04588_),
    .X(_09697_));
 sky130_fd_sc_hd__a21bo_1 _16194_ (.A1(_09693_),
    .A2(_09694_),
    .B1_N(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__nand2_1 _16195_ (.A(_04627_),
    .B(net192),
    .Y(_09699_));
 sky130_fd_sc_hd__nand2_1 _16196_ (.A(_09698_),
    .B(_09699_),
    .Y(_00341_));
 sky130_fd_sc_hd__and3_4 _16197_ (.A(_09554_),
    .B(_09328_),
    .C(_09556_),
    .X(_09700_));
 sky130_fd_sc_hd__clkbuf_2 _16198_ (.A(_09700_),
    .X(_09701_));
 sky130_fd_sc_hd__clkbuf_4 _16199_ (.A(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__mux2_1 _16200_ (.A0(\core.cpuregs[22][0] ),
    .A1(_09315_),
    .S(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__buf_1 _16201_ (.A(_09703_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_4 _16202_ (.A0(\core.cpuregs[22][1] ),
    .A1(_09337_),
    .S(_09702_),
    .X(_09704_));
 sky130_fd_sc_hd__clkbuf_1 _16203_ (.A(_09704_),
    .X(_00343_));
 sky130_fd_sc_hd__clkbuf_2 _16204_ (.A(_09701_),
    .X(_09705_));
 sky130_fd_sc_hd__mux2_1 _16205_ (.A0(\core.cpuregs[22][2] ),
    .A1(_09340_),
    .S(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__buf_1 _16206_ (.A(_09706_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(\core.cpuregs[22][3] ),
    .A1(_09349_),
    .S(_09705_),
    .X(_09707_));
 sky130_fd_sc_hd__buf_1 _16208_ (.A(_09707_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(\core.cpuregs[22][4] ),
    .A1(_09357_),
    .S(_09705_),
    .X(_09708_));
 sky130_fd_sc_hd__clkbuf_1 _16210_ (.A(_09708_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_2 _16211_ (.A0(\core.cpuregs[22][5] ),
    .A1(_09363_),
    .S(_09705_),
    .X(_09709_));
 sky130_fd_sc_hd__buf_1 _16212_ (.A(_09709_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(\core.cpuregs[22][6] ),
    .A1(_09369_),
    .S(_09705_),
    .X(_09710_));
 sky130_fd_sc_hd__clkbuf_1 _16214_ (.A(_09710_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_2 _16215_ (.A0(\core.cpuregs[22][7] ),
    .A1(_09375_),
    .S(_09705_),
    .X(_09711_));
 sky130_fd_sc_hd__clkbuf_1 _16216_ (.A(_09711_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(\core.cpuregs[22][8] ),
    .A1(_09381_),
    .S(_09701_),
    .X(_09712_));
 sky130_fd_sc_hd__buf_1 _16218_ (.A(_09712_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(\core.cpuregs[22][9] ),
    .A1(_09388_),
    .S(_09701_),
    .X(_09713_));
 sky130_fd_sc_hd__clkbuf_2 _16220_ (.A(_09713_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(\core.cpuregs[22][10] ),
    .A1(_09395_),
    .S(_09701_),
    .X(_09714_));
 sky130_fd_sc_hd__buf_1 _16222_ (.A(_09714_),
    .X(_00352_));
 sky130_fd_sc_hd__inv_2 _16223_ (.A(_09700_),
    .Y(_09715_));
 sky130_fd_sc_hd__clkbuf_2 _16224_ (.A(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(_09401_),
    .A1(\core.cpuregs[22][11] ),
    .S(_09716_),
    .X(_09717_));
 sky130_fd_sc_hd__clkbuf_2 _16226_ (.A(_09717_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_8 _16227_ (.A0(\core.cpuregs[22][12] ),
    .A1(_09408_),
    .S(_09701_),
    .X(_09718_));
 sky130_fd_sc_hd__buf_1 _16228_ (.A(_09718_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _16229_ (.A0(_09414_),
    .A1(\core.cpuregs[22][13] ),
    .S(_09716_),
    .X(_09719_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16230_ (.A(_09719_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(_09419_),
    .A1(\core.cpuregs[22][14] ),
    .S(_09715_),
    .X(_09720_));
 sky130_fd_sc_hd__clkbuf_1 _16232_ (.A(_09720_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _16233_ (.A0(_09424_),
    .A1(\core.cpuregs[22][15] ),
    .S(_09715_),
    .X(_09721_));
 sky130_fd_sc_hd__buf_1 _16234_ (.A(_09721_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_8 _16235_ (.A0(_09431_),
    .A1(\core.cpuregs[22][16] ),
    .S(_09715_),
    .X(_09722_));
 sky130_fd_sc_hd__clkbuf_1 _16236_ (.A(_09722_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(_09436_),
    .A1(\core.cpuregs[22][17] ),
    .S(_09715_),
    .X(_09723_));
 sky130_fd_sc_hd__clkbuf_1 _16238_ (.A(_09723_),
    .X(_00359_));
 sky130_fd_sc_hd__nand2_1 _16239_ (.A(_09716_),
    .B(\core.cpuregs[22][18] ),
    .Y(_09724_));
 sky130_fd_sc_hd__a21bo_1 _16240_ (.A1(_09442_),
    .A2(_09702_),
    .B1_N(_09724_),
    .X(_00360_));
 sky130_fd_sc_hd__clkbuf_2 _16241_ (.A(_09702_),
    .X(_09725_));
 sky130_fd_sc_hd__nand2_1 _16242_ (.A(_09448_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__buf_2 _16243_ (.A(_09716_),
    .X(_09727_));
 sky130_fd_sc_hd__nand2_1 _16244_ (.A(_09727_),
    .B(\core.cpuregs[22][19] ),
    .Y(_09728_));
 sky130_fd_sc_hd__nand2_1 _16245_ (.A(_09726_),
    .B(_09728_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_2 _16246_ (.A(_09458_),
    .B(_09725_),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_1 _16247_ (.A(_09727_),
    .B(\core.cpuregs[22][20] ),
    .Y(_09730_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(_09729_),
    .B(_09730_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_2 _16249_ (.A(_09467_),
    .B(_09725_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(_09727_),
    .B(\core.cpuregs[22][21] ),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_1 _16251_ (.A(_09731_),
    .B(_09732_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _16252_ (.A(_09474_),
    .B(_09725_),
    .Y(_09733_));
 sky130_fd_sc_hd__nand2_1 _16253_ (.A(_09727_),
    .B(\core.cpuregs[22][22] ),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _16254_ (.A(_09733_),
    .B(_09734_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _16255_ (.A(_09481_),
    .B(_09725_),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(_09727_),
    .B(\core.cpuregs[22][23] ),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_1 _16257_ (.A(_09735_),
    .B(_09736_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(_09489_),
    .B(_09725_),
    .Y(_09737_));
 sky130_fd_sc_hd__nand2_1 _16259_ (.A(_09727_),
    .B(\core.cpuregs[22][24] ),
    .Y(_09738_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_09737_),
    .B(_09738_),
    .Y(_00366_));
 sky130_fd_sc_hd__clkbuf_4 _16261_ (.A(_09702_),
    .X(_09739_));
 sky130_fd_sc_hd__nand2_1 _16262_ (.A(_09499_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__buf_4 _16263_ (.A(_09716_),
    .X(_09741_));
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(_09741_),
    .B(\core.cpuregs[22][25] ),
    .Y(_09742_));
 sky130_fd_sc_hd__nand2_1 _16265_ (.A(_09740_),
    .B(_09742_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(_09509_),
    .B(_09739_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_2 _16267_ (.A(_09741_),
    .B(\core.cpuregs[22][26] ),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_1 _16268_ (.A(_09743_),
    .B(_09744_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _16269_ (.A(_09516_),
    .B(_09739_),
    .Y(_09745_));
 sky130_fd_sc_hd__nand2_1 _16270_ (.A(_09741_),
    .B(\core.cpuregs[22][27] ),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _16271_ (.A(_09745_),
    .B(_09746_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _16272_ (.A(_09525_),
    .B(_09739_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand2_1 _16273_ (.A(_09741_),
    .B(\core.cpuregs[22][28] ),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_1 _16274_ (.A(_09747_),
    .B(_09748_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_2 _16275_ (.A(_09534_),
    .B(_09739_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(_09741_),
    .B(\core.cpuregs[22][29] ),
    .Y(_09750_));
 sky130_fd_sc_hd__nand2_1 _16277_ (.A(_09749_),
    .B(_09750_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _16278_ (.A(_09542_),
    .B(_09739_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2_1 _16279_ (.A(_09741_),
    .B(\core.cpuregs[22][30] ),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_1 _16280_ (.A(_09751_),
    .B(_09752_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_1 _16281_ (.A(_09551_),
    .B(_09702_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand2_1 _16282_ (.A(_09716_),
    .B(net152),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(_09753_),
    .B(_09754_),
    .Y(_00373_));
 sky130_fd_sc_hd__and3_4 _16284_ (.A(_09554_),
    .B(_09320_),
    .C(_09556_),
    .X(_09755_));
 sky130_fd_sc_hd__clkbuf_2 _16285_ (.A(_09755_),
    .X(_09756_));
 sky130_fd_sc_hd__clkbuf_2 _16286_ (.A(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(\core.cpuregs[2][0] ),
    .A1(_09315_),
    .S(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16288_ (.A(_09758_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_2 _16289_ (.A0(\core.cpuregs[2][1] ),
    .A1(_09337_),
    .S(_09757_),
    .X(_09759_));
 sky130_fd_sc_hd__clkbuf_1 _16290_ (.A(_09759_),
    .X(_00375_));
 sky130_fd_sc_hd__clkbuf_4 _16291_ (.A(_09756_),
    .X(_09760_));
 sky130_fd_sc_hd__mux2_1 _16292_ (.A0(\core.cpuregs[2][2] ),
    .A1(_09340_),
    .S(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__clkbuf_1 _16293_ (.A(_09761_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _16294_ (.A0(\core.cpuregs[2][3] ),
    .A1(_09349_),
    .S(_09760_),
    .X(_09762_));
 sky130_fd_sc_hd__buf_1 _16295_ (.A(_09762_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_2 _16296_ (.A0(\core.cpuregs[2][4] ),
    .A1(_09357_),
    .S(_09760_),
    .X(_09763_));
 sky130_fd_sc_hd__buf_1 _16297_ (.A(_09763_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _16298_ (.A0(\core.cpuregs[2][5] ),
    .A1(_09363_),
    .S(_09760_),
    .X(_09764_));
 sky130_fd_sc_hd__buf_1 _16299_ (.A(_09764_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_2 _16300_ (.A0(\core.cpuregs[2][6] ),
    .A1(_09369_),
    .S(_09760_),
    .X(_09765_));
 sky130_fd_sc_hd__buf_1 _16301_ (.A(_09765_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _16302_ (.A0(\core.cpuregs[2][7] ),
    .A1(_09375_),
    .S(_09760_),
    .X(_09766_));
 sky130_fd_sc_hd__buf_1 _16303_ (.A(_09766_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _16304_ (.A0(\core.cpuregs[2][8] ),
    .A1(_09381_),
    .S(_09756_),
    .X(_09767_));
 sky130_fd_sc_hd__clkbuf_1 _16305_ (.A(_09767_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _16306_ (.A0(\core.cpuregs[2][9] ),
    .A1(_09388_),
    .S(_09756_),
    .X(_09768_));
 sky130_fd_sc_hd__clkbuf_1 _16307_ (.A(_09768_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_4 _16308_ (.A0(\core.cpuregs[2][10] ),
    .A1(_09395_),
    .S(_09756_),
    .X(_09769_));
 sky130_fd_sc_hd__buf_1 _16309_ (.A(_09769_),
    .X(_00384_));
 sky130_fd_sc_hd__inv_2 _16310_ (.A(_09755_),
    .Y(_09770_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16311_ (.A(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__mux2_1 _16312_ (.A0(_09401_),
    .A1(\core.cpuregs[2][11] ),
    .S(_09771_),
    .X(_09772_));
 sky130_fd_sc_hd__clkbuf_1 _16313_ (.A(_09772_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _16314_ (.A0(\core.cpuregs[2][12] ),
    .A1(_09408_),
    .S(_09756_),
    .X(_09773_));
 sky130_fd_sc_hd__buf_1 _16315_ (.A(_09773_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _16316_ (.A0(_09414_),
    .A1(\core.cpuregs[2][13] ),
    .S(_09771_),
    .X(_09774_));
 sky130_fd_sc_hd__clkbuf_1 _16317_ (.A(_09774_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(_09419_),
    .A1(\core.cpuregs[2][14] ),
    .S(_09770_),
    .X(_09775_));
 sky130_fd_sc_hd__clkbuf_1 _16319_ (.A(_09775_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(_09424_),
    .A1(\core.cpuregs[2][15] ),
    .S(_09770_),
    .X(_09776_));
 sky130_fd_sc_hd__clkbuf_1 _16321_ (.A(_09776_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _16322_ (.A0(_09431_),
    .A1(\core.cpuregs[2][16] ),
    .S(_09770_),
    .X(_09777_));
 sky130_fd_sc_hd__clkbuf_1 _16323_ (.A(_09777_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(_09436_),
    .A1(\core.cpuregs[2][17] ),
    .S(_09770_),
    .X(_09778_));
 sky130_fd_sc_hd__clkbuf_1 _16325_ (.A(_09778_),
    .X(_00391_));
 sky130_fd_sc_hd__clkbuf_4 _16326_ (.A(_09441_),
    .X(_09779_));
 sky130_fd_sc_hd__and2_1 _16327_ (.A(_09771_),
    .B(\core.cpuregs[2][18] ),
    .X(_09780_));
 sky130_fd_sc_hd__a21o_1 _16328_ (.A1(_09779_),
    .A2(_09757_),
    .B1(_09780_),
    .X(_00392_));
 sky130_fd_sc_hd__clkbuf_4 _16329_ (.A(_09757_),
    .X(_09781_));
 sky130_fd_sc_hd__nand2_1 _16330_ (.A(_09448_),
    .B(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__clkbuf_4 _16331_ (.A(_09771_),
    .X(_09783_));
 sky130_fd_sc_hd__nand2_1 _16332_ (.A(_09783_),
    .B(net161),
    .Y(_09784_));
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(_09782_),
    .B(_09784_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_2 _16334_ (.A(_09458_),
    .B(_09781_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand2_1 _16335_ (.A(_09783_),
    .B(\core.cpuregs[2][20] ),
    .Y(_09786_));
 sky130_fd_sc_hd__nand2_1 _16336_ (.A(_09785_),
    .B(_09786_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_2 _16337_ (.A(_09467_),
    .B(_09781_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(_09783_),
    .B(net193),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_1 _16339_ (.A(_09787_),
    .B(_09788_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _16340_ (.A(_09474_),
    .B(_09781_),
    .Y(_09789_));
 sky130_fd_sc_hd__nand2_1 _16341_ (.A(_09783_),
    .B(\core.cpuregs[2][22] ),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(_09789_),
    .B(_09790_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(_09481_),
    .B(_09781_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(_09783_),
    .B(net162),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_1 _16345_ (.A(_09791_),
    .B(_09792_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_2 _16346_ (.A(_09489_),
    .B(_09781_),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_1 _16347_ (.A(_09783_),
    .B(\core.cpuregs[2][24] ),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(_09793_),
    .B(_09794_),
    .Y(_00398_));
 sky130_fd_sc_hd__buf_4 _16349_ (.A(_09757_),
    .X(_09795_));
 sky130_fd_sc_hd__nand2_4 _16350_ (.A(_09499_),
    .B(_09795_),
    .Y(_09796_));
 sky130_fd_sc_hd__clkbuf_2 _16351_ (.A(_09771_),
    .X(_09797_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(_09797_),
    .B(net179),
    .Y(_09798_));
 sky130_fd_sc_hd__nand2_1 _16353_ (.A(_09796_),
    .B(_09798_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _16354_ (.A(_09509_),
    .B(_09795_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(_09797_),
    .B(\core.cpuregs[2][26] ),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_1 _16356_ (.A(_09799_),
    .B(_09800_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _16357_ (.A(_09516_),
    .B(_09795_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand2_1 _16358_ (.A(_09797_),
    .B(\core.cpuregs[2][27] ),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_1 _16359_ (.A(_09801_),
    .B(_09802_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_4 _16360_ (.A(_09525_),
    .B(_09795_),
    .Y(_09803_));
 sky130_fd_sc_hd__nand2_1 _16361_ (.A(_09797_),
    .B(\core.cpuregs[2][28] ),
    .Y(_09804_));
 sky130_fd_sc_hd__nand2_1 _16362_ (.A(_09803_),
    .B(_09804_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_4 _16363_ (.A(_09534_),
    .B(_09795_),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_2 _16364_ (.A(_09797_),
    .B(\core.cpuregs[2][29] ),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_2 _16365_ (.A(_09805_),
    .B(_09806_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(_09542_),
    .B(_09795_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand2_2 _16367_ (.A(_09797_),
    .B(\core.cpuregs[2][30] ),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_1 _16368_ (.A(_09807_),
    .B(_09808_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _16369_ (.A(_09551_),
    .B(_09757_),
    .Y(_09809_));
 sky130_fd_sc_hd__nand2_1 _16370_ (.A(_09771_),
    .B(net189),
    .Y(_09810_));
 sky130_fd_sc_hd__nand2_1 _16371_ (.A(_09809_),
    .B(_09810_),
    .Y(_00405_));
 sky130_fd_sc_hd__or3_2 _16372_ (.A(\core.latched_rd[2] ),
    .B(_09317_),
    .C(_09318_),
    .X(_09811_));
 sky130_fd_sc_hd__nand2_4 _16373_ (.A(_09323_),
    .B(_09326_),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_2 _16374_ (.A(_09811_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__clkbuf_2 _16375_ (.A(_09813_),
    .X(_09814_));
 sky130_fd_sc_hd__clkbuf_2 _16376_ (.A(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__mux2_8 _16377_ (.A0(\core.cpuregs[27][0] ),
    .A1(_09315_),
    .S(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__clkbuf_1 _16378_ (.A(_09816_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(\core.cpuregs[27][1] ),
    .A1(_09337_),
    .S(_09815_),
    .X(_09817_));
 sky130_fd_sc_hd__clkbuf_1 _16380_ (.A(_09817_),
    .X(_00407_));
 sky130_fd_sc_hd__clkbuf_4 _16381_ (.A(_09814_),
    .X(_09818_));
 sky130_fd_sc_hd__mux2_1 _16382_ (.A0(\core.cpuregs[27][2] ),
    .A1(_09340_),
    .S(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__buf_1 _16383_ (.A(_09819_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _16384_ (.A0(\core.cpuregs[27][3] ),
    .A1(_09349_),
    .S(_09818_),
    .X(_09820_));
 sky130_fd_sc_hd__buf_1 _16385_ (.A(_09820_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _16386_ (.A0(\core.cpuregs[27][4] ),
    .A1(_09357_),
    .S(_09818_),
    .X(_09821_));
 sky130_fd_sc_hd__buf_1 _16387_ (.A(_09821_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _16388_ (.A0(\core.cpuregs[27][5] ),
    .A1(_09363_),
    .S(_09818_),
    .X(_09822_));
 sky130_fd_sc_hd__clkbuf_1 _16389_ (.A(_09822_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _16390_ (.A0(\core.cpuregs[27][6] ),
    .A1(_09369_),
    .S(_09818_),
    .X(_09823_));
 sky130_fd_sc_hd__buf_1 _16391_ (.A(_09823_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _16392_ (.A0(\core.cpuregs[27][7] ),
    .A1(_09375_),
    .S(_09818_),
    .X(_09824_));
 sky130_fd_sc_hd__clkbuf_1 _16393_ (.A(_09824_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _16394_ (.A0(\core.cpuregs[27][8] ),
    .A1(_09381_),
    .S(_09814_),
    .X(_09825_));
 sky130_fd_sc_hd__clkbuf_1 _16395_ (.A(_09825_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _16396_ (.A0(\core.cpuregs[27][9] ),
    .A1(_09388_),
    .S(_09814_),
    .X(_09826_));
 sky130_fd_sc_hd__buf_1 _16397_ (.A(_09826_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _16398_ (.A0(\core.cpuregs[27][10] ),
    .A1(_09395_),
    .S(_09814_),
    .X(_09827_));
 sky130_fd_sc_hd__clkbuf_1 _16399_ (.A(_09827_),
    .X(_00416_));
 sky130_fd_sc_hd__inv_2 _16400_ (.A(_09813_),
    .Y(_09828_));
 sky130_fd_sc_hd__clkbuf_4 _16401_ (.A(_09828_),
    .X(_09829_));
 sky130_fd_sc_hd__mux2_1 _16402_ (.A0(_09401_),
    .A1(\core.cpuregs[27][11] ),
    .S(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__buf_1 _16403_ (.A(_09830_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_4 _16404_ (.A0(\core.cpuregs[27][12] ),
    .A1(_09408_),
    .S(_09814_),
    .X(_09831_));
 sky130_fd_sc_hd__clkbuf_1 _16405_ (.A(_09831_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _16406_ (.A0(_09414_),
    .A1(\core.cpuregs[27][13] ),
    .S(_09829_),
    .X(_09832_));
 sky130_fd_sc_hd__clkbuf_1 _16407_ (.A(_09832_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(_09419_),
    .A1(\core.cpuregs[27][14] ),
    .S(_09828_),
    .X(_09833_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16409_ (.A(_09833_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_4 _16410_ (.A0(_09424_),
    .A1(\core.cpuregs[27][15] ),
    .S(_09828_),
    .X(_09834_));
 sky130_fd_sc_hd__clkbuf_1 _16411_ (.A(_09834_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _16412_ (.A0(_09431_),
    .A1(\core.cpuregs[27][16] ),
    .S(_09828_),
    .X(_09835_));
 sky130_fd_sc_hd__clkbuf_1 _16413_ (.A(_09835_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_4 _16414_ (.A0(_09436_),
    .A1(\core.cpuregs[27][17] ),
    .S(_09828_),
    .X(_09836_));
 sky130_fd_sc_hd__clkbuf_1 _16415_ (.A(_09836_),
    .X(_00423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16416_ (.A(_09441_),
    .X(_09837_));
 sky130_fd_sc_hd__nand2_4 _16417_ (.A(_09829_),
    .B(\core.cpuregs[27][18] ),
    .Y(_09838_));
 sky130_fd_sc_hd__a21bo_1 _16418_ (.A1(_09837_),
    .A2(_09815_),
    .B1_N(_09838_),
    .X(_00424_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16419_ (.A(_09815_),
    .X(_09839_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(_09448_),
    .B(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16421_ (.A(_09829_),
    .X(_09841_));
 sky130_fd_sc_hd__nand2_1 _16422_ (.A(_09841_),
    .B(net196),
    .Y(_09842_));
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(_09840_),
    .B(_09842_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _16424_ (.A(_09458_),
    .B(_09839_),
    .Y(_09843_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(_09841_),
    .B(net129),
    .Y(_09844_));
 sky130_fd_sc_hd__nand2_1 _16426_ (.A(_09843_),
    .B(_09844_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(_09467_),
    .B(_09839_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_1 _16428_ (.A(_09841_),
    .B(\core.cpuregs[27][21] ),
    .Y(_09846_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(_09845_),
    .B(_09846_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_2 _16430_ (.A(_09474_),
    .B(_09839_),
    .Y(_09847_));
 sky130_fd_sc_hd__nand2_1 _16431_ (.A(_09841_),
    .B(net158),
    .Y(_09848_));
 sky130_fd_sc_hd__nand2_2 _16432_ (.A(_09847_),
    .B(_09848_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_09481_),
    .B(_09839_),
    .Y(_09849_));
 sky130_fd_sc_hd__nand2_1 _16434_ (.A(_09841_),
    .B(net185),
    .Y(_09850_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(_09849_),
    .B(_09850_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _16436_ (.A(_09489_),
    .B(_09839_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand2_1 _16437_ (.A(_09841_),
    .B(\core.cpuregs[27][24] ),
    .Y(_09852_));
 sky130_fd_sc_hd__nand2_1 _16438_ (.A(_09851_),
    .B(_09852_),
    .Y(_00430_));
 sky130_fd_sc_hd__clkbuf_4 _16439_ (.A(_09815_),
    .X(_09853_));
 sky130_fd_sc_hd__nand2_1 _16440_ (.A(_09499_),
    .B(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16441_ (.A(_09829_),
    .X(_09855_));
 sky130_fd_sc_hd__nand2_1 _16442_ (.A(_09855_),
    .B(\core.cpuregs[27][25] ),
    .Y(_09856_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(_09854_),
    .B(_09856_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _16444_ (.A(_09509_),
    .B(_09853_),
    .Y(_09857_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(_09855_),
    .B(\core.cpuregs[27][26] ),
    .Y(_09858_));
 sky130_fd_sc_hd__nand2_1 _16446_ (.A(_09857_),
    .B(_09858_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(_09516_),
    .B(_09853_),
    .Y(_09859_));
 sky130_fd_sc_hd__nand2_1 _16448_ (.A(_09855_),
    .B(\core.cpuregs[27][27] ),
    .Y(_09860_));
 sky130_fd_sc_hd__nand2_1 _16449_ (.A(_09859_),
    .B(_09860_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _16450_ (.A(_09525_),
    .B(_09853_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(_09855_),
    .B(\core.cpuregs[27][28] ),
    .Y(_09862_));
 sky130_fd_sc_hd__nand2_1 _16452_ (.A(_09861_),
    .B(_09862_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(_09534_),
    .B(_09853_),
    .Y(_09863_));
 sky130_fd_sc_hd__nand2_1 _16454_ (.A(_09855_),
    .B(\core.cpuregs[27][29] ),
    .Y(_09864_));
 sky130_fd_sc_hd__nand2_1 _16455_ (.A(_09863_),
    .B(_09864_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_2 _16456_ (.A(_09542_),
    .B(_09853_),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_1 _16457_ (.A(_09855_),
    .B(\core.cpuregs[27][30] ),
    .Y(_09866_));
 sky130_fd_sc_hd__nand2_2 _16458_ (.A(_09865_),
    .B(_09866_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _16459_ (.A(_09551_),
    .B(_09815_),
    .Y(_09867_));
 sky130_fd_sc_hd__nand2_8 _16460_ (.A(_09829_),
    .B(\core.cpuregs[27][31] ),
    .Y(_09868_));
 sky130_fd_sc_hd__nand2_2 _16461_ (.A(_09867_),
    .B(_09868_),
    .Y(_00437_));
 sky130_fd_sc_hd__or3_1 _16462_ (.A(_04370_),
    .B(_04513_),
    .C(_05968_),
    .X(_09869_));
 sky130_fd_sc_hd__nor2_1 _16463_ (.A(_09296_),
    .B(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__clkbuf_2 _16464_ (.A(_09870_),
    .X(_09871_));
 sky130_fd_sc_hd__buf_4 _16465_ (.A(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__mux2_1 _16466_ (.A0(net67),
    .A1(_04694_),
    .S(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__clkbuf_1 _16467_ (.A(_09873_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _16468_ (.A0(net78),
    .A1(_04696_),
    .S(_09872_),
    .X(_09874_));
 sky130_fd_sc_hd__clkbuf_1 _16469_ (.A(_09874_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _16470_ (.A0(net89),
    .A1(\core.mem_la_wdata[2] ),
    .S(_09872_),
    .X(_09875_));
 sky130_fd_sc_hd__clkbuf_1 _16471_ (.A(_09875_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _16472_ (.A0(net92),
    .A1(_04679_),
    .S(_09872_),
    .X(_09876_));
 sky130_fd_sc_hd__clkbuf_1 _16473_ (.A(_09876_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _16474_ (.A0(net93),
    .A1(_04722_),
    .S(_09872_),
    .X(_09877_));
 sky130_fd_sc_hd__clkbuf_1 _16475_ (.A(_09877_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _16476_ (.A0(net94),
    .A1(_04714_),
    .S(_09872_),
    .X(_09878_));
 sky130_fd_sc_hd__clkbuf_1 _16477_ (.A(_09878_),
    .X(_00443_));
 sky130_fd_sc_hd__clkbuf_2 _16478_ (.A(_09871_),
    .X(_09879_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(net95),
    .A1(_04709_),
    .S(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__clkbuf_1 _16480_ (.A(_09880_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _16481_ (.A0(net96),
    .A1(_04705_),
    .S(_09879_),
    .X(_09881_));
 sky130_fd_sc_hd__clkbuf_1 _16482_ (.A(_09881_),
    .X(_00445_));
 sky130_fd_sc_hd__clkbuf_2 _16483_ (.A(_05172_),
    .X(_09882_));
 sky130_fd_sc_hd__clkbuf_2 _16484_ (.A(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__a22o_1 _16485_ (.A1(_04411_),
    .A2(_04694_),
    .B1(_04516_),
    .B2(\core.pcpi_rs2[8] ),
    .X(_09884_));
 sky130_fd_sc_hd__a21o_1 _16486_ (.A1(\core.pcpi_rs2[8] ),
    .A2(_09883_),
    .B1(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(net97),
    .A1(_09885_),
    .S(_09879_),
    .X(_09886_));
 sky130_fd_sc_hd__clkbuf_1 _16488_ (.A(_09886_),
    .X(_00446_));
 sky130_fd_sc_hd__a22o_1 _16489_ (.A1(_04411_),
    .A2(_04696_),
    .B1(_04516_),
    .B2(\core.pcpi_rs2[9] ),
    .X(_09887_));
 sky130_fd_sc_hd__a21o_1 _16490_ (.A1(\core.pcpi_rs2[9] ),
    .A2(_09883_),
    .B1(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(net98),
    .A1(_09888_),
    .S(_09879_),
    .X(_09889_));
 sky130_fd_sc_hd__clkbuf_1 _16492_ (.A(_09889_),
    .X(_00447_));
 sky130_fd_sc_hd__a22o_1 _16493_ (.A1(_04411_),
    .A2(\core.mem_la_wdata[2] ),
    .B1(_04516_),
    .B2(\core.pcpi_rs2[10] ),
    .X(_09890_));
 sky130_fd_sc_hd__a21o_1 _16494_ (.A1(\core.pcpi_rs2[10] ),
    .A2(_09883_),
    .B1(_09890_),
    .X(_09891_));
 sky130_fd_sc_hd__mux2_2 _16495_ (.A0(net68),
    .A1(_09891_),
    .S(_09879_),
    .X(_09892_));
 sky130_fd_sc_hd__clkbuf_1 _16496_ (.A(_09892_),
    .X(_00448_));
 sky130_fd_sc_hd__a22o_1 _16497_ (.A1(_05083_),
    .A2(_04679_),
    .B1(_04516_),
    .B2(\core.pcpi_rs2[11] ),
    .X(_09893_));
 sky130_fd_sc_hd__a21o_1 _16498_ (.A1(\core.pcpi_rs2[11] ),
    .A2(_09883_),
    .B1(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__mux2_1 _16499_ (.A0(net69),
    .A1(_09894_),
    .S(_09879_),
    .X(_09895_));
 sky130_fd_sc_hd__clkbuf_1 _16500_ (.A(_09895_),
    .X(_00449_));
 sky130_fd_sc_hd__a22o_1 _16501_ (.A1(_05083_),
    .A2(_04722_),
    .B1(_04516_),
    .B2(\core.pcpi_rs2[12] ),
    .X(_09896_));
 sky130_fd_sc_hd__a21o_1 _16502_ (.A1(\core.pcpi_rs2[12] ),
    .A2(_09883_),
    .B1(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__buf_4 _16503_ (.A(_09871_),
    .X(_09898_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(net70),
    .A1(_09897_),
    .S(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__buf_1 _16505_ (.A(_09899_),
    .X(_00450_));
 sky130_fd_sc_hd__a22o_2 _16506_ (.A1(_05083_),
    .A2(_04714_),
    .B1(_05174_),
    .B2(\core.pcpi_rs2[13] ),
    .X(_09900_));
 sky130_fd_sc_hd__a21o_1 _16507_ (.A1(\core.pcpi_rs2[13] ),
    .A2(_09883_),
    .B1(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(net71),
    .A1(_09901_),
    .S(_09898_),
    .X(_09902_));
 sky130_fd_sc_hd__clkbuf_1 _16509_ (.A(_09902_),
    .X(_00451_));
 sky130_fd_sc_hd__clkbuf_2 _16510_ (.A(_09882_),
    .X(_09903_));
 sky130_fd_sc_hd__a22o_1 _16511_ (.A1(_05083_),
    .A2(_04709_),
    .B1(_05174_),
    .B2(\core.pcpi_rs2[14] ),
    .X(_09904_));
 sky130_fd_sc_hd__a21o_4 _16512_ (.A1(\core.pcpi_rs2[14] ),
    .A2(_09903_),
    .B1(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__mux2_1 _16513_ (.A0(net72),
    .A1(_09905_),
    .S(_09898_),
    .X(_09906_));
 sky130_fd_sc_hd__clkbuf_1 _16514_ (.A(_09906_),
    .X(_00452_));
 sky130_fd_sc_hd__a22o_1 _16515_ (.A1(_05083_),
    .A2(_04705_),
    .B1(_05174_),
    .B2(\core.pcpi_rs2[15] ),
    .X(_09907_));
 sky130_fd_sc_hd__a21o_1 _16516_ (.A1(\core.pcpi_rs2[15] ),
    .A2(_09903_),
    .B1(_09907_),
    .X(_09908_));
 sky130_fd_sc_hd__mux2_1 _16517_ (.A0(net73),
    .A1(_09908_),
    .S(_09898_),
    .X(_09909_));
 sky130_fd_sc_hd__clkbuf_1 _16518_ (.A(_09909_),
    .X(_00453_));
 sky130_fd_sc_hd__buf_2 _16519_ (.A(_05172_),
    .X(_09910_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(_04694_),
    .A1(\core.pcpi_rs2[16] ),
    .S(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__mux2_1 _16521_ (.A0(net74),
    .A1(_09911_),
    .S(_09898_),
    .X(_09912_));
 sky130_fd_sc_hd__buf_1 _16522_ (.A(_09912_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _16523_ (.A0(_04696_),
    .A1(\core.pcpi_rs2[17] ),
    .S(_09910_),
    .X(_09913_));
 sky130_fd_sc_hd__mux2_1 _16524_ (.A0(net75),
    .A1(_09913_),
    .S(_09898_),
    .X(_09914_));
 sky130_fd_sc_hd__buf_1 _16525_ (.A(_09914_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _16526_ (.A0(\core.mem_la_wdata[2] ),
    .A1(\core.pcpi_rs2[18] ),
    .S(_09910_),
    .X(_09915_));
 sky130_fd_sc_hd__buf_4 _16527_ (.A(_09871_),
    .X(_09916_));
 sky130_fd_sc_hd__mux2_1 _16528_ (.A0(net76),
    .A1(_09915_),
    .S(_09916_),
    .X(_09917_));
 sky130_fd_sc_hd__clkbuf_1 _16529_ (.A(_09917_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _16530_ (.A0(_04679_),
    .A1(\core.pcpi_rs2[19] ),
    .S(_09910_),
    .X(_09918_));
 sky130_fd_sc_hd__mux2_1 _16531_ (.A0(net77),
    .A1(_09918_),
    .S(_09916_),
    .X(_09919_));
 sky130_fd_sc_hd__clkbuf_1 _16532_ (.A(_09919_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _16533_ (.A0(_04722_),
    .A1(\core.pcpi_rs2[20] ),
    .S(_09910_),
    .X(_09920_));
 sky130_fd_sc_hd__mux2_1 _16534_ (.A0(net79),
    .A1(_09920_),
    .S(_09916_),
    .X(_09921_));
 sky130_fd_sc_hd__clkbuf_1 _16535_ (.A(_09921_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _16536_ (.A0(_04714_),
    .A1(\core.pcpi_rs2[21] ),
    .S(_09910_),
    .X(_09922_));
 sky130_fd_sc_hd__mux2_1 _16537_ (.A0(net80),
    .A1(_09922_),
    .S(_09916_),
    .X(_09923_));
 sky130_fd_sc_hd__clkbuf_1 _16538_ (.A(_09923_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _16539_ (.A0(_04709_),
    .A1(\core.pcpi_rs2[22] ),
    .S(_09882_),
    .X(_09924_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(net81),
    .A1(_09924_),
    .S(_09916_),
    .X(_09925_));
 sky130_fd_sc_hd__clkbuf_1 _16541_ (.A(_09925_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _16542_ (.A0(_04705_),
    .A1(\core.pcpi_rs2[23] ),
    .S(_09882_),
    .X(_09926_));
 sky130_fd_sc_hd__mux2_1 _16543_ (.A0(net82),
    .A1(_09926_),
    .S(_09916_),
    .X(_09927_));
 sky130_fd_sc_hd__buf_1 _16544_ (.A(_09927_),
    .X(_00461_));
 sky130_fd_sc_hd__a21o_1 _16545_ (.A1(\core.pcpi_rs2[24] ),
    .A2(_09903_),
    .B1(_09884_),
    .X(_09928_));
 sky130_fd_sc_hd__clkbuf_2 _16546_ (.A(_09870_),
    .X(_09929_));
 sky130_fd_sc_hd__mux2_1 _16547_ (.A0(net83),
    .A1(_09928_),
    .S(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__clkbuf_1 _16548_ (.A(_09930_),
    .X(_00462_));
 sky130_fd_sc_hd__a21o_1 _16549_ (.A1(\core.pcpi_rs2[25] ),
    .A2(_09903_),
    .B1(_09887_),
    .X(_09931_));
 sky130_fd_sc_hd__mux2_1 _16550_ (.A0(net84),
    .A1(_09931_),
    .S(_09929_),
    .X(_09932_));
 sky130_fd_sc_hd__clkbuf_1 _16551_ (.A(_09932_),
    .X(_00463_));
 sky130_fd_sc_hd__a21o_1 _16552_ (.A1(\core.pcpi_rs2[26] ),
    .A2(_09903_),
    .B1(_09890_),
    .X(_09933_));
 sky130_fd_sc_hd__mux2_1 _16553_ (.A0(net85),
    .A1(_09933_),
    .S(_09929_),
    .X(_09934_));
 sky130_fd_sc_hd__clkbuf_1 _16554_ (.A(_09934_),
    .X(_00464_));
 sky130_fd_sc_hd__a21o_1 _16555_ (.A1(\core.pcpi_rs2[27] ),
    .A2(_09903_),
    .B1(_09893_),
    .X(_09935_));
 sky130_fd_sc_hd__mux2_1 _16556_ (.A0(net86),
    .A1(_09935_),
    .S(_09929_),
    .X(_09936_));
 sky130_fd_sc_hd__clkbuf_1 _16557_ (.A(_09936_),
    .X(_00465_));
 sky130_fd_sc_hd__a21o_1 _16558_ (.A1(\core.pcpi_rs2[28] ),
    .A2(_05424_),
    .B1(_09896_),
    .X(_09937_));
 sky130_fd_sc_hd__mux2_1 _16559_ (.A0(net87),
    .A1(_09937_),
    .S(_09929_),
    .X(_09938_));
 sky130_fd_sc_hd__clkbuf_1 _16560_ (.A(_09938_),
    .X(_00466_));
 sky130_fd_sc_hd__a21o_1 _16561_ (.A1(\core.pcpi_rs2[29] ),
    .A2(_05424_),
    .B1(_09900_),
    .X(_09939_));
 sky130_fd_sc_hd__mux2_1 _16562_ (.A0(net88),
    .A1(_09939_),
    .S(_09929_),
    .X(_09940_));
 sky130_fd_sc_hd__buf_1 _16563_ (.A(_09940_),
    .X(_00467_));
 sky130_fd_sc_hd__a21o_1 _16564_ (.A1(\core.pcpi_rs2[30] ),
    .A2(_05424_),
    .B1(_09904_),
    .X(_09941_));
 sky130_fd_sc_hd__mux2_1 _16565_ (.A0(net90),
    .A1(_09941_),
    .S(_09871_),
    .X(_09942_));
 sky130_fd_sc_hd__buf_1 _16566_ (.A(_09942_),
    .X(_00468_));
 sky130_fd_sc_hd__a21o_1 _16567_ (.A1(\core.pcpi_rs2[31] ),
    .A2(_05424_),
    .B1(_09907_),
    .X(_09943_));
 sky130_fd_sc_hd__mux2_1 _16568_ (.A0(net91),
    .A1(_09943_),
    .S(_09871_),
    .X(_09944_));
 sky130_fd_sc_hd__clkbuf_1 _16569_ (.A(_09944_),
    .X(_00469_));
 sky130_fd_sc_hd__clkbuf_2 _16570_ (.A(_05972_),
    .X(_09945_));
 sky130_fd_sc_hd__inv_2 _16571_ (.A(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__and3_1 _16572_ (.A(_09946_),
    .B(_04370_),
    .C(_06021_),
    .X(_09947_));
 sky130_fd_sc_hd__a21o_1 _16573_ (.A1(net115),
    .A2(_05973_),
    .B1(_09947_),
    .X(_00470_));
 sky130_fd_sc_hd__inv_2 _16574_ (.A(_09557_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(_09323_),
    .B(_09321_),
    .Y(_09949_));
 sky130_fd_sc_hd__clkbuf_4 _16576_ (.A(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__nor2_1 _16577_ (.A(_09948_),
    .B(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__clkbuf_2 _16578_ (.A(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__clkbuf_2 _16579_ (.A(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__mux2_4 _16580_ (.A0(\core.cpuregs[28][0] ),
    .A1(_09315_),
    .S(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__clkbuf_1 _16581_ (.A(_09954_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _16582_ (.A0(\core.cpuregs[28][1] ),
    .A1(_09337_),
    .S(_09953_),
    .X(_09955_));
 sky130_fd_sc_hd__buf_1 _16583_ (.A(_09955_),
    .X(_00472_));
 sky130_fd_sc_hd__clkbuf_4 _16584_ (.A(_09952_),
    .X(_09956_));
 sky130_fd_sc_hd__mux2_1 _16585_ (.A0(\core.cpuregs[28][2] ),
    .A1(_09340_),
    .S(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__buf_1 _16586_ (.A(_09957_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _16587_ (.A0(\core.cpuregs[28][3] ),
    .A1(_09349_),
    .S(_09956_),
    .X(_09958_));
 sky130_fd_sc_hd__clkbuf_1 _16588_ (.A(_09958_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _16589_ (.A0(\core.cpuregs[28][4] ),
    .A1(_09357_),
    .S(_09956_),
    .X(_09959_));
 sky130_fd_sc_hd__clkbuf_1 _16590_ (.A(_09959_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _16591_ (.A0(\core.cpuregs[28][5] ),
    .A1(_09363_),
    .S(_09956_),
    .X(_09960_));
 sky130_fd_sc_hd__clkbuf_1 _16592_ (.A(_09960_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _16593_ (.A0(\core.cpuregs[28][6] ),
    .A1(_09369_),
    .S(_09956_),
    .X(_09961_));
 sky130_fd_sc_hd__buf_1 _16594_ (.A(_09961_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _16595_ (.A0(\core.cpuregs[28][7] ),
    .A1(_09375_),
    .S(_09956_),
    .X(_09962_));
 sky130_fd_sc_hd__clkbuf_1 _16596_ (.A(_09962_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _16597_ (.A0(\core.cpuregs[28][8] ),
    .A1(_09381_),
    .S(_09952_),
    .X(_09963_));
 sky130_fd_sc_hd__buf_1 _16598_ (.A(_09963_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(\core.cpuregs[28][9] ),
    .A1(_09388_),
    .S(_09952_),
    .X(_09964_));
 sky130_fd_sc_hd__buf_1 _16600_ (.A(_09964_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_2 _16601_ (.A0(\core.cpuregs[28][10] ),
    .A1(_09395_),
    .S(_09952_),
    .X(_09965_));
 sky130_fd_sc_hd__clkbuf_1 _16602_ (.A(_09965_),
    .X(_00481_));
 sky130_fd_sc_hd__inv_2 _16603_ (.A(_09951_),
    .Y(_09966_));
 sky130_fd_sc_hd__buf_2 _16604_ (.A(_09966_),
    .X(_09967_));
 sky130_fd_sc_hd__mux2_1 _16605_ (.A0(_09401_),
    .A1(\core.cpuregs[28][11] ),
    .S(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__clkbuf_1 _16606_ (.A(_09968_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _16607_ (.A0(\core.cpuregs[28][12] ),
    .A1(_09408_),
    .S(_09952_),
    .X(_09969_));
 sky130_fd_sc_hd__buf_1 _16608_ (.A(_09969_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _16609_ (.A0(_09414_),
    .A1(\core.cpuregs[28][13] ),
    .S(_09967_),
    .X(_09970_));
 sky130_fd_sc_hd__buf_1 _16610_ (.A(_09970_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _16611_ (.A0(_09419_),
    .A1(\core.cpuregs[28][14] ),
    .S(_09966_),
    .X(_09971_));
 sky130_fd_sc_hd__clkbuf_1 _16612_ (.A(_09971_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_4 _16613_ (.A0(_09424_),
    .A1(\core.cpuregs[28][15] ),
    .S(_09966_),
    .X(_09972_));
 sky130_fd_sc_hd__clkbuf_1 _16614_ (.A(_09972_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _16615_ (.A0(_09431_),
    .A1(\core.cpuregs[28][16] ),
    .S(_09966_),
    .X(_09973_));
 sky130_fd_sc_hd__buf_1 _16616_ (.A(_09973_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _16617_ (.A0(_09436_),
    .A1(\core.cpuregs[28][17] ),
    .S(_09966_),
    .X(_09974_));
 sky130_fd_sc_hd__clkbuf_1 _16618_ (.A(_09974_),
    .X(_00488_));
 sky130_fd_sc_hd__nand2_8 _16619_ (.A(_09967_),
    .B(\core.cpuregs[28][18] ),
    .Y(_09975_));
 sky130_fd_sc_hd__a21bo_1 _16620_ (.A1(_09837_),
    .A2(_09953_),
    .B1_N(_09975_),
    .X(_00489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16621_ (.A(_09953_),
    .X(_09976_));
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(_09448_),
    .B(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16623_ (.A(_09967_),
    .X(_09978_));
 sky130_fd_sc_hd__nand2_1 _16624_ (.A(_09978_),
    .B(net198),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_1 _16625_ (.A(_09977_),
    .B(_09979_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _16626_ (.A(_09458_),
    .B(_09976_),
    .Y(_09980_));
 sky130_fd_sc_hd__nand2_1 _16627_ (.A(_09978_),
    .B(net124),
    .Y(_09981_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(_09980_),
    .B(_09981_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _16629_ (.A(_09467_),
    .B(_09976_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_1 _16630_ (.A(_09978_),
    .B(\core.cpuregs[28][21] ),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_1 _16631_ (.A(_09982_),
    .B(_09983_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _16632_ (.A(_09474_),
    .B(_09976_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_1 _16633_ (.A(_09978_),
    .B(\core.cpuregs[28][22] ),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2_1 _16634_ (.A(_09984_),
    .B(_09985_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _16635_ (.A(_09481_),
    .B(_09976_),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_1 _16636_ (.A(_09978_),
    .B(\core.cpuregs[28][23] ),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_09986_),
    .B(_09987_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _16638_ (.A(_09489_),
    .B(_09976_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(_09978_),
    .B(\core.cpuregs[28][24] ),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(_09988_),
    .B(_09989_),
    .Y(_00495_));
 sky130_fd_sc_hd__clkbuf_4 _16641_ (.A(_09953_),
    .X(_09990_));
 sky130_fd_sc_hd__nand2_1 _16642_ (.A(_09499_),
    .B(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__clkbuf_2 _16643_ (.A(_09967_),
    .X(_09992_));
 sky130_fd_sc_hd__nand2_2 _16644_ (.A(_09992_),
    .B(\core.cpuregs[28][25] ),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_2 _16645_ (.A(_09991_),
    .B(_09993_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _16646_ (.A(_09509_),
    .B(_09990_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_2 _16647_ (.A(_09992_),
    .B(\core.cpuregs[28][26] ),
    .Y(_09995_));
 sky130_fd_sc_hd__nand2_1 _16648_ (.A(_09994_),
    .B(_09995_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _16649_ (.A(_09516_),
    .B(_09990_),
    .Y(_09996_));
 sky130_fd_sc_hd__nand2_1 _16650_ (.A(_09992_),
    .B(\core.cpuregs[28][27] ),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_1 _16651_ (.A(_09996_),
    .B(_09997_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _16652_ (.A(_09525_),
    .B(_09990_),
    .Y(_09998_));
 sky130_fd_sc_hd__nand2_1 _16653_ (.A(_09992_),
    .B(\core.cpuregs[28][28] ),
    .Y(_09999_));
 sky130_fd_sc_hd__nand2_1 _16654_ (.A(_09998_),
    .B(_09999_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _16655_ (.A(_09534_),
    .B(_09990_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand2_2 _16656_ (.A(_09992_),
    .B(net153),
    .Y(_10001_));
 sky130_fd_sc_hd__nand2_1 _16657_ (.A(_10000_),
    .B(_10001_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(_09542_),
    .B(_09990_),
    .Y(_10002_));
 sky130_fd_sc_hd__nand2_2 _16659_ (.A(_09992_),
    .B(\core.cpuregs[28][30] ),
    .Y(_10003_));
 sky130_fd_sc_hd__nand2_1 _16660_ (.A(_10002_),
    .B(_10003_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _16661_ (.A(_09551_),
    .B(_09953_),
    .Y(_10004_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(_09967_),
    .B(net175),
    .Y(_10005_));
 sky130_fd_sc_hd__nand2_1 _16663_ (.A(_10004_),
    .B(_10005_),
    .Y(_00502_));
 sky130_fd_sc_hd__or2b_1 _16664_ (.A(\core.mem_rdata_q[6] ),
    .B_N(_05939_),
    .X(_10006_));
 sky130_fd_sc_hd__o21a_1 _16665_ (.A1(net29),
    .A2(_05923_),
    .B1(_10006_),
    .X(_10007_));
 sky130_fd_sc_hd__clkbuf_2 _16666_ (.A(_10007_),
    .X(_01349_));
 sky130_fd_sc_hd__inv_2 _16667_ (.A(net27),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_1 _16668_ (.A(_05939_),
    .B(\core.mem_rdata_q[4] ),
    .Y(_10009_));
 sky130_fd_sc_hd__o21ai_1 _16669_ (.A1(_10008_),
    .A2(_05939_),
    .B1(_10009_),
    .Y(_01347_));
 sky130_fd_sc_hd__inv_2 _16670_ (.A(_01347_),
    .Y(_10010_));
 sky130_fd_sc_hd__or2b_1 _16671_ (.A(\core.mem_rdata_q[5] ),
    .B_N(_05922_),
    .X(_10011_));
 sky130_fd_sc_hd__o21a_1 _16672_ (.A1(net28),
    .A2(_05939_),
    .B1(_10011_),
    .X(_10012_));
 sky130_fd_sc_hd__buf_2 _16673_ (.A(_10012_),
    .X(_01348_));
 sky130_fd_sc_hd__inv_2 _16674_ (.A(_01348_),
    .Y(_10013_));
 sky130_fd_sc_hd__or3_1 _16675_ (.A(_01349_),
    .B(_10010_),
    .C(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__inv_2 _16676_ (.A(\core.mem_rdata_q[2] ),
    .Y(_10015_));
 sky130_fd_sc_hd__nand2_1 _16677_ (.A(_05939_),
    .B(_10015_),
    .Y(_10016_));
 sky130_fd_sc_hd__o21a_1 _16678_ (.A1(net23),
    .A2(_05923_),
    .B1(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__buf_4 _16679_ (.A(_10017_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _16680_ (.A0(net26),
    .A1(\core.mem_rdata_q[3] ),
    .S(_05922_),
    .X(_10018_));
 sky130_fd_sc_hd__clkbuf_1 _16681_ (.A(_10018_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _16682_ (.A0(net12),
    .A1(\core.mem_rdata_q[1] ),
    .S(_05922_),
    .X(_10019_));
 sky130_fd_sc_hd__clkbuf_1 _16683_ (.A(_10019_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _16684_ (.A0(net1),
    .A1(\core.mem_rdata_q[0] ),
    .S(_05922_),
    .X(_10020_));
 sky130_fd_sc_hd__clkbuf_1 _16685_ (.A(_10020_),
    .X(_01343_));
 sky130_fd_sc_hd__and2_1 _16686_ (.A(_01344_),
    .B(_01343_),
    .X(_10021_));
 sky130_fd_sc_hd__or2b_1 _16687_ (.A(_01346_),
    .B_N(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__nor2_1 _16688_ (.A(_01345_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__inv_2 _16689_ (.A(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__nor2_1 _16690_ (.A(_10014_),
    .B(_10024_),
    .Y(_10025_));
 sky130_fd_sc_hd__mux2_1 _16691_ (.A0(_10025_),
    .A1(\core.is_alu_reg_reg ),
    .S(_05949_),
    .X(_10026_));
 sky130_fd_sc_hd__clkbuf_1 _16692_ (.A(_10026_),
    .X(_00503_));
 sky130_fd_sc_hd__or3_2 _16693_ (.A(_10010_),
    .B(_01348_),
    .C(_01349_),
    .X(_10027_));
 sky130_fd_sc_hd__nor2_2 _16694_ (.A(_10027_),
    .B(_10024_),
    .Y(_10028_));
 sky130_fd_sc_hd__mux2_2 _16695_ (.A0(_10028_),
    .A1(\core.is_alu_reg_imm ),
    .S(_05949_),
    .X(_10029_));
 sky130_fd_sc_hd__clkbuf_1 _16696_ (.A(_10029_),
    .X(_00504_));
 sky130_fd_sc_hd__inv_2 _16697_ (.A(_01345_),
    .Y(_10030_));
 sky130_fd_sc_hd__nor2_1 _16698_ (.A(_10030_),
    .B(_10022_),
    .Y(_10031_));
 sky130_fd_sc_hd__inv_2 _16699_ (.A(_10031_),
    .Y(_10032_));
 sky130_fd_sc_hd__nor2_1 _16700_ (.A(_10027_),
    .B(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__mux2_1 _16701_ (.A0(_10033_),
    .A1(\core.instr_auipc ),
    .S(_05949_),
    .X(_10034_));
 sky130_fd_sc_hd__clkbuf_1 _16702_ (.A(_10034_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_1 _16703_ (.A(_10014_),
    .B(_10032_),
    .Y(_10035_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(_10035_),
    .A1(_07729_),
    .S(_05949_),
    .X(_10036_));
 sky130_fd_sc_hd__clkbuf_1 _16705_ (.A(_10036_),
    .X(_00506_));
 sky130_fd_sc_hd__o211ai_4 _16706_ (.A1(_04399_),
    .A2(_04380_),
    .B1(_04394_),
    .C1(_04400_),
    .Y(_10037_));
 sky130_fd_sc_hd__or3b_1 _16707_ (.A(_05316_),
    .B(_10037_),
    .C_N(\core.instr_lb ),
    .X(_10038_));
 sky130_fd_sc_hd__nand2_1 _16708_ (.A(_10037_),
    .B(\core.latched_is_lb ),
    .Y(_10039_));
 sky130_fd_sc_hd__a21oi_1 _16709_ (.A1(_10038_),
    .A2(_10039_),
    .B1(_07650_),
    .Y(_00507_));
 sky130_fd_sc_hd__or3_1 _16710_ (.A(_05316_),
    .B(_04426_),
    .C(_10037_),
    .X(_10040_));
 sky130_fd_sc_hd__nand2_1 _16711_ (.A(_10037_),
    .B(\core.latched_is_lh ),
    .Y(_10041_));
 sky130_fd_sc_hd__a21oi_1 _16712_ (.A1(_10040_),
    .A2(_10041_),
    .B1(_07650_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand3_1 _16713_ (.A(_04971_),
    .B(_04975_),
    .C(_04973_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand2_2 _16714_ (.A(_04489_),
    .B(_04425_),
    .Y(_10043_));
 sky130_fd_sc_hd__nand3_1 _16715_ (.A(_10042_),
    .B(_04981_),
    .C(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__buf_1 _16716_ (.A(_04492_),
    .X(_10045_));
 sky130_fd_sc_hd__nand2_2 _16717_ (.A(_06609_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__nand2_4 _16718_ (.A(_10044_),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand2_2 _16719_ (.A(_04492_),
    .B(_04500_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand2_1 _16720_ (.A(_10047_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__or2_1 _16721_ (.A(_09316_),
    .B(_10048_),
    .X(_10050_));
 sky130_fd_sc_hd__a21oi_1 _16722_ (.A1(_10049_),
    .A2(_10050_),
    .B1(_07650_),
    .Y(_00510_));
 sky130_fd_sc_hd__o21ai_1 _16723_ (.A1(_04511_),
    .A2(_04500_),
    .B1(_06601_),
    .Y(_10051_));
 sky130_fd_sc_hd__inv_2 _16724_ (.A(_04505_),
    .Y(_10052_));
 sky130_fd_sc_hd__a21oi_1 _16725_ (.A1(_10051_),
    .A2(_10052_),
    .B1(_07650_),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _16726_ (.A(_04452_),
    .Y(_00512_));
 sky130_fd_sc_hd__nor2_1 _16727_ (.A(\core.decoder_pseudo_trigger ),
    .B(_04501_),
    .Y(_10053_));
 sky130_fd_sc_hd__buf_1 _16728_ (.A(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16729_ (.A(_10054_),
    .X(_10055_));
 sky130_fd_sc_hd__nand2_2 _16730_ (.A(_10054_),
    .B(_04975_),
    .Y(_10056_));
 sky130_fd_sc_hd__inv_2 _16731_ (.A(\core.mem_rdata_q[13] ),
    .Y(_10057_));
 sky130_fd_sc_hd__nand2_2 _16732_ (.A(_10057_),
    .B(\core.mem_rdata_q[12] ),
    .Y(_10058_));
 sky130_fd_sc_hd__nor2_2 _16733_ (.A(\core.mem_rdata_q[14] ),
    .B(_10058_),
    .Y(_10059_));
 sky130_fd_sc_hd__inv_2 _16734_ (.A(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__o22a_1 _16735_ (.A1(_04436_),
    .A2(_10055_),
    .B1(_10056_),
    .B2(_10060_),
    .X(_10061_));
 sky130_fd_sc_hd__nor2_1 _16736_ (.A(_06327_),
    .B(_10061_),
    .Y(_00513_));
 sky130_fd_sc_hd__buf_1 _16737_ (.A(_09314_),
    .X(_10062_));
 sky130_fd_sc_hd__nand2_1 _16738_ (.A(_09555_),
    .B(\core.latched_rd[0] ),
    .Y(_10063_));
 sky130_fd_sc_hd__inv_2 _16739_ (.A(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__and3_1 _16740_ (.A(_09554_),
    .B(_09328_),
    .C(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__clkbuf_2 _16741_ (.A(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__clkbuf_2 _16742_ (.A(_10066_),
    .X(_10067_));
 sky130_fd_sc_hd__mux2_2 _16743_ (.A0(\core.cpuregs[21][0] ),
    .A1(_10062_),
    .S(_10067_),
    .X(_10068_));
 sky130_fd_sc_hd__clkbuf_1 _16744_ (.A(_10068_),
    .X(_00514_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16745_ (.A(_09336_),
    .X(_10069_));
 sky130_fd_sc_hd__mux2_8 _16746_ (.A0(\core.cpuregs[21][1] ),
    .A1(_10069_),
    .S(_10067_),
    .X(_10070_));
 sky130_fd_sc_hd__clkbuf_1 _16747_ (.A(_10070_),
    .X(_00515_));
 sky130_fd_sc_hd__buf_2 _16748_ (.A(_09339_),
    .X(_10071_));
 sky130_fd_sc_hd__clkbuf_2 _16749_ (.A(_10066_),
    .X(_10072_));
 sky130_fd_sc_hd__mux2_1 _16750_ (.A0(\core.cpuregs[21][2] ),
    .A1(_10071_),
    .S(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__buf_1 _16751_ (.A(_10073_),
    .X(_00516_));
 sky130_fd_sc_hd__clkbuf_2 _16752_ (.A(_09348_),
    .X(_10074_));
 sky130_fd_sc_hd__mux2_1 _16753_ (.A0(\core.cpuregs[21][3] ),
    .A1(_10074_),
    .S(_10072_),
    .X(_10075_));
 sky130_fd_sc_hd__buf_1 _16754_ (.A(_10075_),
    .X(_00517_));
 sky130_fd_sc_hd__buf_1 _16755_ (.A(_09356_),
    .X(_10076_));
 sky130_fd_sc_hd__mux2_1 _16756_ (.A0(\core.cpuregs[21][4] ),
    .A1(_10076_),
    .S(_10072_),
    .X(_10077_));
 sky130_fd_sc_hd__clkbuf_1 _16757_ (.A(_10077_),
    .X(_00518_));
 sky130_fd_sc_hd__buf_2 _16758_ (.A(_09362_),
    .X(_10078_));
 sky130_fd_sc_hd__mux2_1 _16759_ (.A0(\core.cpuregs[21][5] ),
    .A1(_10078_),
    .S(_10072_),
    .X(_10079_));
 sky130_fd_sc_hd__clkbuf_1 _16760_ (.A(_10079_),
    .X(_00519_));
 sky130_fd_sc_hd__buf_2 _16761_ (.A(_09368_),
    .X(_10080_));
 sky130_fd_sc_hd__mux2_1 _16762_ (.A0(\core.cpuregs[21][6] ),
    .A1(_10080_),
    .S(_10072_),
    .X(_10081_));
 sky130_fd_sc_hd__clkbuf_1 _16763_ (.A(_10081_),
    .X(_00520_));
 sky130_fd_sc_hd__buf_2 _16764_ (.A(_09374_),
    .X(_10082_));
 sky130_fd_sc_hd__mux2_1 _16765_ (.A0(\core.cpuregs[21][7] ),
    .A1(_10082_),
    .S(_10072_),
    .X(_10083_));
 sky130_fd_sc_hd__clkbuf_1 _16766_ (.A(_10083_),
    .X(_00521_));
 sky130_fd_sc_hd__buf_1 _16767_ (.A(_09380_),
    .X(_10084_));
 sky130_fd_sc_hd__mux2_1 _16768_ (.A0(\core.cpuregs[21][8] ),
    .A1(_10084_),
    .S(_10066_),
    .X(_10085_));
 sky130_fd_sc_hd__clkbuf_1 _16769_ (.A(_10085_),
    .X(_00522_));
 sky130_fd_sc_hd__clkbuf_4 _16770_ (.A(_09387_),
    .X(_10086_));
 sky130_fd_sc_hd__mux2_1 _16771_ (.A0(\core.cpuregs[21][9] ),
    .A1(_10086_),
    .S(_10066_),
    .X(_10087_));
 sky130_fd_sc_hd__buf_1 _16772_ (.A(_10087_),
    .X(_00523_));
 sky130_fd_sc_hd__buf_1 _16773_ (.A(_09394_),
    .X(_10088_));
 sky130_fd_sc_hd__mux2_1 _16774_ (.A0(\core.cpuregs[21][10] ),
    .A1(_10088_),
    .S(_10066_),
    .X(_10089_));
 sky130_fd_sc_hd__clkbuf_1 _16775_ (.A(_10089_),
    .X(_00524_));
 sky130_fd_sc_hd__buf_1 _16776_ (.A(_09400_),
    .X(_10090_));
 sky130_fd_sc_hd__inv_2 _16777_ (.A(_10065_),
    .Y(_10091_));
 sky130_fd_sc_hd__clkbuf_2 _16778_ (.A(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__mux2_2 _16779_ (.A0(_10090_),
    .A1(\core.cpuregs[21][11] ),
    .S(_10092_),
    .X(_10093_));
 sky130_fd_sc_hd__clkbuf_1 _16780_ (.A(_10093_),
    .X(_00525_));
 sky130_fd_sc_hd__buf_1 _16781_ (.A(_09407_),
    .X(_10094_));
 sky130_fd_sc_hd__mux2_2 _16782_ (.A0(\core.cpuregs[21][12] ),
    .A1(_10094_),
    .S(_10066_),
    .X(_10095_));
 sky130_fd_sc_hd__clkbuf_2 _16783_ (.A(_10095_),
    .X(_00526_));
 sky130_fd_sc_hd__buf_1 _16784_ (.A(_09413_),
    .X(_10096_));
 sky130_fd_sc_hd__mux2_1 _16785_ (.A0(_10096_),
    .A1(\core.cpuregs[21][13] ),
    .S(_10092_),
    .X(_10097_));
 sky130_fd_sc_hd__clkbuf_1 _16786_ (.A(_10097_),
    .X(_00527_));
 sky130_fd_sc_hd__buf_1 _16787_ (.A(_09418_),
    .X(_10098_));
 sky130_fd_sc_hd__mux2_4 _16788_ (.A0(_10098_),
    .A1(\core.cpuregs[21][14] ),
    .S(_10091_),
    .X(_10099_));
 sky130_fd_sc_hd__clkbuf_1 _16789_ (.A(_10099_),
    .X(_00528_));
 sky130_fd_sc_hd__buf_1 _16790_ (.A(_09423_),
    .X(_10100_));
 sky130_fd_sc_hd__mux2_4 _16791_ (.A0(_10100_),
    .A1(\core.cpuregs[21][15] ),
    .S(_10091_),
    .X(_10101_));
 sky130_fd_sc_hd__clkbuf_1 _16792_ (.A(_10101_),
    .X(_00529_));
 sky130_fd_sc_hd__buf_1 _16793_ (.A(_09430_),
    .X(_10102_));
 sky130_fd_sc_hd__mux2_1 _16794_ (.A0(_10102_),
    .A1(\core.cpuregs[21][16] ),
    .S(_10091_),
    .X(_10103_));
 sky130_fd_sc_hd__buf_1 _16795_ (.A(_10103_),
    .X(_00530_));
 sky130_fd_sc_hd__clkbuf_4 _16796_ (.A(_09435_),
    .X(_10104_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(_10104_),
    .A1(\core.cpuregs[21][17] ),
    .S(_10091_),
    .X(_10105_));
 sky130_fd_sc_hd__clkbuf_2 _16798_ (.A(_10105_),
    .X(_00531_));
 sky130_fd_sc_hd__nand2_1 _16799_ (.A(_10092_),
    .B(\core.cpuregs[21][18] ),
    .Y(_10106_));
 sky130_fd_sc_hd__a21bo_1 _16800_ (.A1(_09837_),
    .A2(_10067_),
    .B1_N(_10106_),
    .X(_00532_));
 sky130_fd_sc_hd__clkbuf_2 _16801_ (.A(_09447_),
    .X(_10107_));
 sky130_fd_sc_hd__clkbuf_4 _16802_ (.A(_10067_),
    .X(_10108_));
 sky130_fd_sc_hd__nand2_2 _16803_ (.A(_10107_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__clkbuf_4 _16804_ (.A(_10092_),
    .X(_10110_));
 sky130_fd_sc_hd__nand2_1 _16805_ (.A(_10110_),
    .B(\core.cpuregs[21][19] ),
    .Y(_10111_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(_10109_),
    .B(_10111_),
    .Y(_00533_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16807_ (.A(_09457_),
    .X(_10112_));
 sky130_fd_sc_hd__nand2_1 _16808_ (.A(_10112_),
    .B(_10108_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand2_2 _16809_ (.A(_10110_),
    .B(\core.cpuregs[21][20] ),
    .Y(_10114_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(_10113_),
    .B(_10114_),
    .Y(_00534_));
 sky130_fd_sc_hd__buf_6 _16811_ (.A(_09466_),
    .X(_10115_));
 sky130_fd_sc_hd__nand2_1 _16812_ (.A(_10115_),
    .B(_10108_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(_10110_),
    .B(\core.cpuregs[21][21] ),
    .Y(_10117_));
 sky130_fd_sc_hd__nand2_1 _16814_ (.A(_10116_),
    .B(_10117_),
    .Y(_00535_));
 sky130_fd_sc_hd__clkbuf_4 _16815_ (.A(_09473_),
    .X(_10118_));
 sky130_fd_sc_hd__nand2_1 _16816_ (.A(_10118_),
    .B(_10108_),
    .Y(_10119_));
 sky130_fd_sc_hd__nand2_1 _16817_ (.A(_10110_),
    .B(\core.cpuregs[21][22] ),
    .Y(_10120_));
 sky130_fd_sc_hd__nand2_2 _16818_ (.A(_10119_),
    .B(_10120_),
    .Y(_00536_));
 sky130_fd_sc_hd__buf_6 _16819_ (.A(_09480_),
    .X(_10121_));
 sky130_fd_sc_hd__nand2_1 _16820_ (.A(_10121_),
    .B(_10108_),
    .Y(_10122_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(_10110_),
    .B(\core.cpuregs[21][23] ),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_1 _16822_ (.A(_10122_),
    .B(_10123_),
    .Y(_00537_));
 sky130_fd_sc_hd__buf_6 _16823_ (.A(_09488_),
    .X(_10124_));
 sky130_fd_sc_hd__nand2_1 _16824_ (.A(_10124_),
    .B(_10108_),
    .Y(_10125_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(_10110_),
    .B(\core.cpuregs[21][24] ),
    .Y(_10126_));
 sky130_fd_sc_hd__nand2_1 _16826_ (.A(_10125_),
    .B(_10126_),
    .Y(_00538_));
 sky130_fd_sc_hd__buf_2 _16827_ (.A(_09498_),
    .X(_10127_));
 sky130_fd_sc_hd__clkbuf_4 _16828_ (.A(_10067_),
    .X(_10128_));
 sky130_fd_sc_hd__nand2_2 _16829_ (.A(_10127_),
    .B(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__clkbuf_4 _16830_ (.A(_10092_),
    .X(_10130_));
 sky130_fd_sc_hd__nand2_1 _16831_ (.A(_10130_),
    .B(\core.cpuregs[21][25] ),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(_10129_),
    .B(_10131_),
    .Y(_00539_));
 sky130_fd_sc_hd__clkbuf_4 _16833_ (.A(_09508_),
    .X(_10132_));
 sky130_fd_sc_hd__nand2_2 _16834_ (.A(_10132_),
    .B(_10128_),
    .Y(_10133_));
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(_10130_),
    .B(\core.cpuregs[21][26] ),
    .Y(_10134_));
 sky130_fd_sc_hd__nand2_1 _16836_ (.A(_10133_),
    .B(_10134_),
    .Y(_00540_));
 sky130_fd_sc_hd__buf_6 _16837_ (.A(_09515_),
    .X(_10135_));
 sky130_fd_sc_hd__nand2_1 _16838_ (.A(_10135_),
    .B(_10128_),
    .Y(_10136_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(_10130_),
    .B(\core.cpuregs[21][27] ),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_1 _16840_ (.A(_10136_),
    .B(_10137_),
    .Y(_00541_));
 sky130_fd_sc_hd__buf_6 _16841_ (.A(_09524_),
    .X(_10138_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(_10138_),
    .B(_10128_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand2_2 _16843_ (.A(_10130_),
    .B(\core.cpuregs[21][28] ),
    .Y(_10140_));
 sky130_fd_sc_hd__nand2_1 _16844_ (.A(_10139_),
    .B(_10140_),
    .Y(_00542_));
 sky130_fd_sc_hd__clkbuf_4 _16845_ (.A(_09533_),
    .X(_10141_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(_10141_),
    .B(_10128_),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_1 _16847_ (.A(_10130_),
    .B(\core.cpuregs[21][29] ),
    .Y(_10143_));
 sky130_fd_sc_hd__nand2_1 _16848_ (.A(_10142_),
    .B(_10143_),
    .Y(_00543_));
 sky130_fd_sc_hd__buf_6 _16849_ (.A(_09541_),
    .X(_10144_));
 sky130_fd_sc_hd__nand2_2 _16850_ (.A(_10144_),
    .B(_10128_),
    .Y(_10145_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(_10130_),
    .B(net190),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_1 _16852_ (.A(_10145_),
    .B(_10146_),
    .Y(_00544_));
 sky130_fd_sc_hd__clkbuf_2 _16853_ (.A(_09550_),
    .X(_10147_));
 sky130_fd_sc_hd__nand2_1 _16854_ (.A(_10147_),
    .B(_10067_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand2_1 _16855_ (.A(_10092_),
    .B(\core.cpuregs[21][31] ),
    .Y(_10149_));
 sky130_fd_sc_hd__nand2_1 _16856_ (.A(_10148_),
    .B(_10149_),
    .Y(_00545_));
 sky130_fd_sc_hd__and3_1 _16857_ (.A(_01348_),
    .B(_01349_),
    .C(_10010_),
    .X(_10150_));
 sky130_fd_sc_hd__and4_1 _16858_ (.A(_10150_),
    .B(_10021_),
    .C(_01345_),
    .D(_01346_),
    .X(_10151_));
 sky130_fd_sc_hd__mux2_1 _16859_ (.A0(_10151_),
    .A1(_06974_),
    .S(_05949_),
    .X(_10152_));
 sky130_fd_sc_hd__clkbuf_1 _16860_ (.A(_10152_),
    .X(_00546_));
 sky130_fd_sc_hd__inv_2 _16861_ (.A(\core.mem_rdata_q[12] ),
    .Y(_10153_));
 sky130_fd_sc_hd__inv_2 _16862_ (.A(\core.mem_rdata_q[14] ),
    .Y(_10154_));
 sky130_fd_sc_hd__and3_2 _16863_ (.A(_10153_),
    .B(_10057_),
    .C(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__inv_2 _16864_ (.A(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__o22a_1 _16865_ (.A1(_04423_),
    .A2(_10055_),
    .B1(_10056_),
    .B2(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__nor2_2 _16866_ (.A(_06327_),
    .B(_10157_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(_09324_),
    .B(_09556_),
    .Y(_10158_));
 sky130_fd_sc_hd__nor2_1 _16868_ (.A(_09811_),
    .B(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__clkbuf_2 _16869_ (.A(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__clkbuf_2 _16870_ (.A(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__mux2_2 _16871_ (.A0(\core.cpuregs[26][0] ),
    .A1(_10062_),
    .S(_10161_),
    .X(_10162_));
 sky130_fd_sc_hd__clkbuf_1 _16872_ (.A(_10162_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_4 _16873_ (.A0(\core.cpuregs[26][1] ),
    .A1(_10069_),
    .S(_10161_),
    .X(_10163_));
 sky130_fd_sc_hd__clkbuf_1 _16874_ (.A(_10163_),
    .X(_00549_));
 sky130_fd_sc_hd__clkbuf_2 _16875_ (.A(_10160_),
    .X(_10164_));
 sky130_fd_sc_hd__mux2_1 _16876_ (.A0(\core.cpuregs[26][2] ),
    .A1(_10071_),
    .S(_10164_),
    .X(_10165_));
 sky130_fd_sc_hd__buf_1 _16877_ (.A(_10165_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _16878_ (.A0(\core.cpuregs[26][3] ),
    .A1(_10074_),
    .S(_10164_),
    .X(_10166_));
 sky130_fd_sc_hd__buf_1 _16879_ (.A(_10166_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_2 _16880_ (.A0(\core.cpuregs[26][4] ),
    .A1(_10076_),
    .S(_10164_),
    .X(_10167_));
 sky130_fd_sc_hd__buf_1 _16881_ (.A(_10167_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(\core.cpuregs[26][5] ),
    .A1(_10078_),
    .S(_10164_),
    .X(_10168_));
 sky130_fd_sc_hd__clkbuf_1 _16883_ (.A(_10168_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _16884_ (.A0(\core.cpuregs[26][6] ),
    .A1(_10080_),
    .S(_10164_),
    .X(_10169_));
 sky130_fd_sc_hd__clkbuf_1 _16885_ (.A(_10169_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _16886_ (.A0(\core.cpuregs[26][7] ),
    .A1(_10082_),
    .S(_10164_),
    .X(_10170_));
 sky130_fd_sc_hd__buf_1 _16887_ (.A(_10170_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _16888_ (.A0(\core.cpuregs[26][8] ),
    .A1(_10084_),
    .S(_10160_),
    .X(_10171_));
 sky130_fd_sc_hd__clkbuf_1 _16889_ (.A(_10171_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_2 _16890_ (.A0(\core.cpuregs[26][9] ),
    .A1(_10086_),
    .S(_10160_),
    .X(_10172_));
 sky130_fd_sc_hd__buf_1 _16891_ (.A(_10172_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _16892_ (.A0(\core.cpuregs[26][10] ),
    .A1(_10088_),
    .S(_10160_),
    .X(_10173_));
 sky130_fd_sc_hd__clkbuf_1 _16893_ (.A(_10173_),
    .X(_00558_));
 sky130_fd_sc_hd__clkinv_4 _16894_ (.A(_10159_),
    .Y(_10174_));
 sky130_fd_sc_hd__clkbuf_2 _16895_ (.A(_10174_),
    .X(_10175_));
 sky130_fd_sc_hd__mux2_1 _16896_ (.A0(_10090_),
    .A1(\core.cpuregs[26][11] ),
    .S(_10175_),
    .X(_10176_));
 sky130_fd_sc_hd__buf_1 _16897_ (.A(_10176_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_4 _16898_ (.A0(\core.cpuregs[26][12] ),
    .A1(_10094_),
    .S(_10160_),
    .X(_10177_));
 sky130_fd_sc_hd__clkbuf_1 _16899_ (.A(_10177_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _16900_ (.A0(_10096_),
    .A1(\core.cpuregs[26][13] ),
    .S(_10175_),
    .X(_10178_));
 sky130_fd_sc_hd__clkbuf_1 _16901_ (.A(_10178_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _16902_ (.A0(_10098_),
    .A1(\core.cpuregs[26][14] ),
    .S(_10174_),
    .X(_10179_));
 sky130_fd_sc_hd__clkbuf_1 _16903_ (.A(_10179_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_4 _16904_ (.A0(_10100_),
    .A1(\core.cpuregs[26][15] ),
    .S(_10174_),
    .X(_10180_));
 sky130_fd_sc_hd__buf_1 _16905_ (.A(_10180_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _16906_ (.A0(_10102_),
    .A1(\core.cpuregs[26][16] ),
    .S(_10174_),
    .X(_10181_));
 sky130_fd_sc_hd__clkbuf_1 _16907_ (.A(_10181_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_2 _16908_ (.A0(_10104_),
    .A1(\core.cpuregs[26][17] ),
    .S(_10174_),
    .X(_10182_));
 sky130_fd_sc_hd__clkbuf_1 _16909_ (.A(_10182_),
    .X(_00565_));
 sky130_fd_sc_hd__nand2_1 _16910_ (.A(_10175_),
    .B(\core.cpuregs[26][18] ),
    .Y(_10183_));
 sky130_fd_sc_hd__a21bo_1 _16911_ (.A1(_09837_),
    .A2(_10161_),
    .B1_N(_10183_),
    .X(_00566_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16912_ (.A(_10161_),
    .X(_10184_));
 sky130_fd_sc_hd__nand2_1 _16913_ (.A(_10107_),
    .B(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__clkbuf_2 _16914_ (.A(_10175_),
    .X(_10186_));
 sky130_fd_sc_hd__nand2_1 _16915_ (.A(_10186_),
    .B(\core.cpuregs[26][19] ),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_1 _16916_ (.A(_10185_),
    .B(_10187_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(_10112_),
    .B(_10184_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand2_1 _16918_ (.A(_10186_),
    .B(\core.cpuregs[26][20] ),
    .Y(_10189_));
 sky130_fd_sc_hd__nand2_1 _16919_ (.A(_10188_),
    .B(_10189_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _16920_ (.A(_10115_),
    .B(_10184_),
    .Y(_10190_));
 sky130_fd_sc_hd__nand2_4 _16921_ (.A(_10186_),
    .B(\core.cpuregs[26][21] ),
    .Y(_10191_));
 sky130_fd_sc_hd__nand2_1 _16922_ (.A(_10190_),
    .B(_10191_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _16923_ (.A(_10118_),
    .B(_10184_),
    .Y(_10192_));
 sky130_fd_sc_hd__nand2_1 _16924_ (.A(_10186_),
    .B(\core.cpuregs[26][22] ),
    .Y(_10193_));
 sky130_fd_sc_hd__nand2_1 _16925_ (.A(_10192_),
    .B(_10193_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _16926_ (.A(_10121_),
    .B(_10184_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand2_1 _16927_ (.A(_10186_),
    .B(\core.cpuregs[26][23] ),
    .Y(_10195_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(_10194_),
    .B(_10195_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _16929_ (.A(_10124_),
    .B(_10184_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(_10186_),
    .B(\core.cpuregs[26][24] ),
    .Y(_10197_));
 sky130_fd_sc_hd__nand2_1 _16931_ (.A(_10196_),
    .B(_10197_),
    .Y(_00572_));
 sky130_fd_sc_hd__clkbuf_4 _16932_ (.A(_10161_),
    .X(_10198_));
 sky130_fd_sc_hd__nand2_1 _16933_ (.A(_10127_),
    .B(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__clkbuf_2 _16934_ (.A(_10175_),
    .X(_10200_));
 sky130_fd_sc_hd__nand2_1 _16935_ (.A(_10200_),
    .B(\core.cpuregs[26][25] ),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(_10199_),
    .B(_10201_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _16937_ (.A(_10132_),
    .B(_10198_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(_10200_),
    .B(\core.cpuregs[26][26] ),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_1 _16939_ (.A(_10202_),
    .B(_10203_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(_10135_),
    .B(_10198_),
    .Y(_10204_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_10200_),
    .B(\core.cpuregs[26][27] ),
    .Y(_10205_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(_10204_),
    .B(_10205_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_2 _16943_ (.A(_10138_),
    .B(_10198_),
    .Y(_10206_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(_10200_),
    .B(\core.cpuregs[26][28] ),
    .Y(_10207_));
 sky130_fd_sc_hd__nand2_1 _16945_ (.A(_10206_),
    .B(_10207_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(_10141_),
    .B(_10198_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_4 _16947_ (.A(_10200_),
    .B(\core.cpuregs[26][29] ),
    .Y(_10209_));
 sky130_fd_sc_hd__nand2_1 _16948_ (.A(_10208_),
    .B(_10209_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _16949_ (.A(_10144_),
    .B(_10198_),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_2 _16950_ (.A(_10200_),
    .B(\core.cpuregs[26][30] ),
    .Y(_10211_));
 sky130_fd_sc_hd__nand2_1 _16951_ (.A(_10210_),
    .B(_10211_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _16952_ (.A(_10147_),
    .B(_10161_),
    .Y(_10212_));
 sky130_fd_sc_hd__nand2_1 _16953_ (.A(_10175_),
    .B(\core.cpuregs[26][31] ),
    .Y(_10213_));
 sky130_fd_sc_hd__nand2_1 _16954_ (.A(_10212_),
    .B(_10213_),
    .Y(_00579_));
 sky130_fd_sc_hd__inv_2 _16955_ (.A(_10053_),
    .Y(_10214_));
 sky130_fd_sc_hd__buf_1 _16956_ (.A(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__buf_2 _16957_ (.A(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__buf_1 _16958_ (.A(_10216_),
    .X(_10217_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _16959_ (.A(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(_10054_),
    .B(_04468_),
    .Y(_10219_));
 sky130_fd_sc_hd__inv_2 _16961_ (.A(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__a22o_1 _16962_ (.A1(\core.instr_sh ),
    .A2(_10218_),
    .B1(_10220_),
    .B2(_10059_),
    .X(_00580_));
 sky130_fd_sc_hd__nand2_2 _16963_ (.A(_10053_),
    .B(\core.is_alu_reg_imm ),
    .Y(_10221_));
 sky130_fd_sc_hd__and3_1 _16964_ (.A(_10153_),
    .B(_10154_),
    .C(\core.mem_rdata_q[13] ),
    .X(_10222_));
 sky130_fd_sc_hd__inv_2 _16965_ (.A(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__o22a_1 _16966_ (.A1(_04422_),
    .A2(_10055_),
    .B1(_10221_),
    .B2(_10223_),
    .X(_10224_));
 sky130_fd_sc_hd__nor2_1 _16967_ (.A(_06327_),
    .B(_10224_),
    .Y(_00581_));
 sky130_fd_sc_hd__clkbuf_2 _16968_ (.A(_10214_),
    .X(_10225_));
 sky130_fd_sc_hd__clkbuf_2 _16969_ (.A(_10225_),
    .X(_10226_));
 sky130_fd_sc_hd__or3_1 _16970_ (.A(\core.mem_rdata_q[14] ),
    .B(_10153_),
    .C(_10057_),
    .X(_10227_));
 sky130_fd_sc_hd__o2bb2a_1 _16971_ (.A1_N(\core.instr_sltiu ),
    .A2_N(_10226_),
    .B1(_10221_),
    .B2(_10227_),
    .X(_10228_));
 sky130_fd_sc_hd__nor2_1 _16972_ (.A(_06327_),
    .B(_10228_),
    .Y(_00582_));
 sky130_fd_sc_hd__or3_1 _16973_ (.A(\core.mem_rdata_q[12] ),
    .B(_10057_),
    .C(_10154_),
    .X(_10229_));
 sky130_fd_sc_hd__o2bb2a_1 _16974_ (.A1_N(\core.instr_ori ),
    .A2_N(_10226_),
    .B1(_10221_),
    .B2(_10229_),
    .X(_10230_));
 sky130_fd_sc_hd__nor2_1 _16975_ (.A(_06327_),
    .B(_10230_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(_10042_),
    .B(_05194_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand3_1 _16977_ (.A(_10231_),
    .B(_05068_),
    .C(_06314_),
    .Y(_10232_));
 sky130_fd_sc_hd__nor2_1 _16978_ (.A(_04391_),
    .B(\core.cpu_state[2] ),
    .Y(_10233_));
 sky130_fd_sc_hd__a22o_1 _16979_ (.A1(_04992_),
    .A2(_10233_),
    .B1(_04465_),
    .B2(_04466_),
    .X(_10234_));
 sky130_fd_sc_hd__inv_2 _16980_ (.A(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand2_1 _16981_ (.A(_10232_),
    .B(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_2 _16982_ (.A(_10234_),
    .B(\core.latched_store ),
    .Y(_10237_));
 sky130_fd_sc_hd__a21oi_1 _16983_ (.A1(_10236_),
    .A2(_10237_),
    .B1(_07650_),
    .Y(_00584_));
 sky130_fd_sc_hd__clkbuf_2 _16984_ (.A(\core.mem_rdata_q[31] ),
    .X(_10238_));
 sky130_fd_sc_hd__nor2_1 _16985_ (.A(\core.mem_rdata_q[26] ),
    .B(\core.mem_rdata_q[27] ),
    .Y(_10239_));
 sky130_fd_sc_hd__inv_2 _16986_ (.A(\core.mem_rdata_q[25] ),
    .Y(_10240_));
 sky130_fd_sc_hd__inv_2 _16987_ (.A(\core.mem_rdata_q[28] ),
    .Y(_10241_));
 sky130_fd_sc_hd__and3_1 _16988_ (.A(_10239_),
    .B(_10240_),
    .C(_10241_),
    .X(_10242_));
 sky130_fd_sc_hd__inv_2 _16989_ (.A(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__or4_2 _16990_ (.A(\core.mem_rdata_q[29] ),
    .B(\core.mem_rdata_q[30] ),
    .C(_10238_),
    .D(_10243_),
    .X(_10244_));
 sky130_fd_sc_hd__clkbuf_2 _16991_ (.A(_10244_),
    .X(_10245_));
 sky130_fd_sc_hd__inv_2 _16992_ (.A(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__buf_2 _16993_ (.A(_10054_),
    .X(_10247_));
 sky130_fd_sc_hd__or2_2 _16994_ (.A(_10154_),
    .B(_10058_),
    .X(_10248_));
 sky130_fd_sc_hd__inv_2 _16995_ (.A(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__and2_1 _16996_ (.A(_10249_),
    .B(\core.is_alu_reg_imm ),
    .X(_10250_));
 sky130_fd_sc_hd__and2_1 _16997_ (.A(_10217_),
    .B(\core.instr_srli ),
    .X(_10251_));
 sky130_fd_sc_hd__a31o_1 _16998_ (.A1(_10246_),
    .A2(_10247_),
    .A3(_10250_),
    .B1(_10251_),
    .X(_00585_));
 sky130_fd_sc_hd__nand2_1 _16999_ (.A(_10155_),
    .B(\core.is_alu_reg_reg ),
    .Y(_10252_));
 sky130_fd_sc_hd__or3_1 _17000_ (.A(_10225_),
    .B(_10252_),
    .C(_10245_),
    .X(_10253_));
 sky130_fd_sc_hd__buf_2 _17001_ (.A(_10216_),
    .X(_10254_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(_10254_),
    .B(\core.instr_add ),
    .Y(_10255_));
 sky130_fd_sc_hd__clkbuf_2 _17003_ (.A(_04514_),
    .X(_10256_));
 sky130_fd_sc_hd__a21oi_1 _17004_ (.A1(_10253_),
    .A2(_10255_),
    .B1(_10256_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_2 _17005_ (.A(_10053_),
    .B(\core.is_alu_reg_reg ),
    .Y(_10257_));
 sky130_fd_sc_hd__or3_1 _17006_ (.A(_10060_),
    .B(_10257_),
    .C(_10245_),
    .X(_10258_));
 sky130_fd_sc_hd__nand2_1 _17007_ (.A(_10254_),
    .B(\core.instr_sll ),
    .Y(_10259_));
 sky130_fd_sc_hd__a21oi_1 _17008_ (.A1(_10258_),
    .A2(_10259_),
    .B1(_10256_),
    .Y(_00587_));
 sky130_fd_sc_hd__and3_1 _17009_ (.A(_10153_),
    .B(_10057_),
    .C(\core.mem_rdata_q[14] ),
    .X(_10260_));
 sky130_fd_sc_hd__inv_2 _17010_ (.A(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__or3_1 _17011_ (.A(_10257_),
    .B(_10261_),
    .C(_10245_),
    .X(_10262_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(_10254_),
    .B(\core.instr_xor ),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_1 _17013_ (.A1(_10262_),
    .A2(_10263_),
    .B1(_10256_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(_10249_),
    .B(\core.is_alu_reg_reg ),
    .Y(_10264_));
 sky130_fd_sc_hd__inv_2 _17015_ (.A(\core.mem_rdata_q[31] ),
    .Y(_10265_));
 sky130_fd_sc_hd__inv_2 _17016_ (.A(\core.mem_rdata_q[30] ),
    .Y(_10266_));
 sky130_fd_sc_hd__nor2_1 _17017_ (.A(\core.mem_rdata_q[29] ),
    .B(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__and3_2 _17018_ (.A(_10242_),
    .B(_10265_),
    .C(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__inv_2 _17019_ (.A(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__or3_1 _17020_ (.A(_10225_),
    .B(_10264_),
    .C(_10269_),
    .X(_10270_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(_10254_),
    .B(\core.instr_sra ),
    .Y(_10271_));
 sky130_fd_sc_hd__a21oi_1 _17022_ (.A1(_10270_),
    .A2(_10271_),
    .B1(_10256_),
    .Y(_00589_));
 sky130_fd_sc_hd__nor2_1 _17023_ (.A(_04975_),
    .B(\core.instr_sltiu ),
    .Y(_10272_));
 sky130_fd_sc_hd__a311o_2 _17024_ (.A1(_04414_),
    .A2(_10272_),
    .A3(_04422_),
    .B1(_06325_),
    .C1(_10055_),
    .X(_10273_));
 sky130_fd_sc_hd__inv_2 _17025_ (.A(_10273_),
    .Y(_00590_));
 sky130_fd_sc_hd__and2_1 _17026_ (.A(_10045_),
    .B(\core.decoded_rd[0] ),
    .X(_10274_));
 sky130_fd_sc_hd__and3_4 _17027_ (.A(_10052_),
    .B(_04388_),
    .C(_10048_),
    .X(_10275_));
 sky130_fd_sc_hd__mux2_4 _17028_ (.A0(\core.latched_rd[0] ),
    .A1(_10274_),
    .S(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__clkbuf_2 _17029_ (.A(_10276_),
    .X(_00591_));
 sky130_fd_sc_hd__and2_1 _17030_ (.A(_10045_),
    .B(\core.decoded_rd[1] ),
    .X(_10277_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(\core.latched_rd[1] ),
    .A1(_10277_),
    .S(_10275_),
    .X(_10278_));
 sky130_fd_sc_hd__clkbuf_1 _17032_ (.A(_10278_),
    .X(_00592_));
 sky130_fd_sc_hd__and2_1 _17033_ (.A(_10045_),
    .B(\core.decoded_rd[2] ),
    .X(_10279_));
 sky130_fd_sc_hd__mux2_4 _17034_ (.A0(\core.latched_rd[2] ),
    .A1(_10279_),
    .S(_10275_),
    .X(_10280_));
 sky130_fd_sc_hd__clkbuf_1 _17035_ (.A(_10280_),
    .X(_00593_));
 sky130_fd_sc_hd__and2_1 _17036_ (.A(_10045_),
    .B(\core.decoded_rd[3] ),
    .X(_10281_));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(\core.latched_rd[3] ),
    .A1(_10281_),
    .S(_10275_),
    .X(_10282_));
 sky130_fd_sc_hd__clkbuf_1 _17038_ (.A(_10282_),
    .X(_00594_));
 sky130_fd_sc_hd__and2_1 _17039_ (.A(_10045_),
    .B(\core.decoded_rd[4] ),
    .X(_10283_));
 sky130_fd_sc_hd__mux2_4 _17040_ (.A0(\core.latched_rd[4] ),
    .A1(_10283_),
    .S(_10275_),
    .X(_10284_));
 sky130_fd_sc_hd__clkbuf_1 _17041_ (.A(_10284_),
    .X(_00595_));
 sky130_fd_sc_hd__inv_2 _17042_ (.A(_09869_),
    .Y(_10285_));
 sky130_fd_sc_hd__o21a_1 _17043_ (.A1(_05968_),
    .A2(_05967_),
    .B1(_09295_),
    .X(_10286_));
 sky130_fd_sc_hd__a32o_1 _17044_ (.A1(_05029_),
    .A2(_10285_),
    .A3(_10286_),
    .B1(_05973_),
    .B2(net118),
    .X(_00596_));
 sky130_fd_sc_hd__o21ai_2 _17045_ (.A1(_04693_),
    .A2(_05047_),
    .B1(_04996_),
    .Y(_10287_));
 sky130_fd_sc_hd__a32o_1 _17046_ (.A1(_10285_),
    .A2(_10286_),
    .A3(_10287_),
    .B1(_05973_),
    .B2(net109),
    .X(_00597_));
 sky130_fd_sc_hd__or3_1 _17047_ (.A(_09882_),
    .B(_05028_),
    .C(_05033_),
    .X(_10288_));
 sky130_fd_sc_hd__a32o_1 _17048_ (.A1(_10285_),
    .A2(_10286_),
    .A3(_10288_),
    .B1(_05973_),
    .B2(net101),
    .X(_00598_));
 sky130_fd_sc_hd__or3_1 _17049_ (.A(_09882_),
    .B(_05005_),
    .C(_05028_),
    .X(_10289_));
 sky130_fd_sc_hd__a32o_1 _17050_ (.A1(_10285_),
    .A2(_10286_),
    .A3(_10289_),
    .B1(_05973_),
    .B2(net114),
    .X(_00599_));
 sky130_fd_sc_hd__or3_1 _17051_ (.A(\core.mem_rdata_q[17] ),
    .B(\core.mem_rdata_q[18] ),
    .C(\core.mem_rdata_q[19] ),
    .X(_10290_));
 sky130_fd_sc_hd__or3_1 _17052_ (.A(\core.mem_rdata_q[15] ),
    .B(\core.mem_rdata_q[16] ),
    .C(_10290_),
    .X(_10291_));
 sky130_fd_sc_hd__nor2_1 _17053_ (.A(_10223_),
    .B(_10291_),
    .Y(_10292_));
 sky130_fd_sc_hd__inv_2 _17054_ (.A(\core.mem_rdata_q[24] ),
    .Y(_10293_));
 sky130_fd_sc_hd__inv_2 _17055_ (.A(\core.mem_rdata_q[27] ),
    .Y(_10294_));
 sky130_fd_sc_hd__nor2_4 _17056_ (.A(\core.mem_rdata_q[26] ),
    .B(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__and4_1 _17057_ (.A(_10292_),
    .B(_10293_),
    .C(_10240_),
    .D(_10295_),
    .X(_10296_));
 sky130_fd_sc_hd__nand2_1 _17058_ (.A(\core.mem_rdata_q[0] ),
    .B(\core.mem_rdata_q[1] ),
    .Y(_10297_));
 sky130_fd_sc_hd__inv_2 _17059_ (.A(\core.mem_rdata_q[3] ),
    .Y(_10298_));
 sky130_fd_sc_hd__and4_1 _17060_ (.A(_10241_),
    .B(_10015_),
    .C(_10298_),
    .D(_10238_),
    .X(_10299_));
 sky130_fd_sc_hd__and3_1 _17061_ (.A(\core.mem_rdata_q[4] ),
    .B(\core.mem_rdata_q[5] ),
    .C(\core.mem_rdata_q[6] ),
    .X(_10300_));
 sky130_fd_sc_hd__and4b_1 _17062_ (.A_N(_10297_),
    .B(_10299_),
    .C(_10267_),
    .D(_10300_),
    .X(_10301_));
 sky130_fd_sc_hd__inv_2 _17063_ (.A(\core.mem_rdata_q[21] ),
    .Y(_10302_));
 sky130_fd_sc_hd__inv_2 _17064_ (.A(\core.mem_rdata_q[22] ),
    .Y(_10303_));
 sky130_fd_sc_hd__inv_2 _17065_ (.A(\core.mem_rdata_q[23] ),
    .Y(_10304_));
 sky130_fd_sc_hd__and4_1 _17066_ (.A(_10054_),
    .B(_10302_),
    .C(_10303_),
    .D(_10304_),
    .X(_10305_));
 sky130_fd_sc_hd__clkbuf_2 _17067_ (.A(_10217_),
    .X(_10306_));
 sky130_fd_sc_hd__a32o_1 _17068_ (.A1(_10296_),
    .A2(_10301_),
    .A3(_10305_),
    .B1(_05142_),
    .B2(_10306_),
    .X(_00600_));
 sky130_fd_sc_hd__o32a_1 _17069_ (.A1(_04374_),
    .A2(_04375_),
    .A3(_09297_),
    .B1(net33),
    .B2(_09302_),
    .X(_10307_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(_09301_),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__a21o_1 _17071_ (.A1(_10308_),
    .A2(net66),
    .B1(_09946_),
    .X(_00601_));
 sky130_fd_sc_hd__or3_1 _17072_ (.A(\core.mem_rdata_q[4] ),
    .B(\core.mem_rdata_q[5] ),
    .C(\core.mem_rdata_q[6] ),
    .X(_10309_));
 sky130_fd_sc_hd__or3_1 _17073_ (.A(_10015_),
    .B(_10298_),
    .C(_10297_),
    .X(_10310_));
 sky130_fd_sc_hd__or4_1 _17074_ (.A(_10225_),
    .B(_10156_),
    .C(_10309_),
    .D(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__buf_2 _17075_ (.A(_10216_),
    .X(_10312_));
 sky130_fd_sc_hd__nand2_1 _17076_ (.A(_10312_),
    .B(\core.instr_fence ),
    .Y(_10313_));
 sky130_fd_sc_hd__a21oi_1 _17077_ (.A1(_10311_),
    .A2(_10313_),
    .B1(_10256_),
    .Y(_00602_));
 sky130_fd_sc_hd__and2b_1 _17078_ (.A_N(\core.cpu_state[0] ),
    .B(_06614_),
    .X(_10314_));
 sky130_fd_sc_hd__nand3_1 _17079_ (.A(_04993_),
    .B(_10314_),
    .C(_04439_),
    .Y(_10315_));
 sky130_fd_sc_hd__or2_2 _17080_ (.A(_04513_),
    .B(_04377_),
    .X(_10316_));
 sky130_fd_sc_hd__inv_2 _17081_ (.A(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__a2bb2o_1 _17082_ (.A1_N(_10315_),
    .A2_N(_04381_),
    .B1(\core.mem_do_wdata ),
    .B2(_10317_),
    .X(_00603_));
 sky130_fd_sc_hd__buf_2 _17083_ (.A(_04496_),
    .X(_10318_));
 sky130_fd_sc_hd__nand2_1 _17084_ (.A(_10318_),
    .B(\core.decoded_imm[0] ),
    .Y(_10319_));
 sky130_fd_sc_hd__o21ai_1 _17085_ (.A1(_04498_),
    .A2(_09655_),
    .B1(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__nand2_1 _17086_ (.A(_04387_),
    .B(\core.cpu_state[2] ),
    .Y(_10321_));
 sky130_fd_sc_hd__clkbuf_4 _17087_ (.A(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__mux2_1 _17088_ (.A0(_10320_),
    .A1(_04694_),
    .S(_10322_),
    .X(_10323_));
 sky130_fd_sc_hd__clkbuf_1 _17089_ (.A(_10323_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _17090_ (.A(_10318_),
    .B(\core.decoded_imm[1] ),
    .Y(_10324_));
 sky130_fd_sc_hd__o21ai_2 _17091_ (.A1(_04498_),
    .A2(_09692_),
    .B1(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__mux2_1 _17092_ (.A0(_10325_),
    .A1(_04696_),
    .S(_10322_),
    .X(_10326_));
 sky130_fd_sc_hd__clkbuf_1 _17093_ (.A(_10326_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _17094_ (.A(_10318_),
    .B(\core.decoded_imm[2] ),
    .Y(_10327_));
 sky130_fd_sc_hd__o21ai_2 _17095_ (.A1(_04498_),
    .A2(_04583_),
    .B1(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__mux2_1 _17096_ (.A0(_10328_),
    .A1(\core.mem_la_wdata[2] ),
    .S(_10322_),
    .X(_10329_));
 sky130_fd_sc_hd__buf_4 _17097_ (.A(_10329_),
    .X(_00606_));
 sky130_fd_sc_hd__nand2_1 _17098_ (.A(_10318_),
    .B(\core.decoded_imm[3] ),
    .Y(_10330_));
 sky130_fd_sc_hd__o21ai_2 _17099_ (.A1(_04498_),
    .A2(_04623_),
    .B1(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__mux2_1 _17100_ (.A0(_10331_),
    .A1(_04679_),
    .S(_10322_),
    .X(_10332_));
 sky130_fd_sc_hd__clkbuf_4 _17101_ (.A(_10332_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _17102_ (.A(_10318_),
    .B(\core.decoded_imm[4] ),
    .Y(_10333_));
 sky130_fd_sc_hd__o21ai_1 _17103_ (.A1(_04498_),
    .A2(_04675_),
    .B1(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__mux2_1 _17104_ (.A0(_10334_),
    .A1(_04722_),
    .S(_10322_),
    .X(_10335_));
 sky130_fd_sc_hd__buf_4 _17105_ (.A(_10335_),
    .X(_00608_));
 sky130_fd_sc_hd__buf_1 _17106_ (.A(_00004_),
    .X(_10336_));
 sky130_fd_sc_hd__buf_2 _17107_ (.A(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17108_ (.A(_04520_),
    .X(_10338_));
 sky130_fd_sc_hd__clkbuf_2 _17109_ (.A(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__clkbuf_2 _17110_ (.A(_10339_),
    .X(_10340_));
 sky130_fd_sc_hd__mux2_1 _17111_ (.A0(\core.cpuregs[24][5] ),
    .A1(\core.cpuregs[25][5] ),
    .S(_10340_),
    .X(_10341_));
 sky130_fd_sc_hd__clkbuf_2 _17112_ (.A(_04567_),
    .X(_10342_));
 sky130_fd_sc_hd__mux2_1 _17113_ (.A0(\core.cpuregs[26][5] ),
    .A1(\core.cpuregs[27][5] ),
    .S(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__clkbuf_2 _17114_ (.A(_04641_),
    .X(_10344_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(_10341_),
    .A1(_10343_),
    .S(_10344_),
    .X(_10345_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17116_ (.A(_04549_),
    .X(_10346_));
 sky130_fd_sc_hd__clkbuf_8 _17117_ (.A(_10346_),
    .X(_10347_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17118_ (.A(_10347_),
    .X(_10348_));
 sky130_fd_sc_hd__nand2_1 _17119_ (.A(_10345_),
    .B(_10348_),
    .Y(_10349_));
 sky130_fd_sc_hd__clkbuf_2 _17120_ (.A(_04662_),
    .X(_10350_));
 sky130_fd_sc_hd__mux2_1 _17121_ (.A0(\core.cpuregs[28][5] ),
    .A1(\core.cpuregs[29][5] ),
    .S(_10350_),
    .X(_10351_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17122_ (.A(_04531_),
    .X(_10352_));
 sky130_fd_sc_hd__clkbuf_2 _17123_ (.A(_10352_),
    .X(_10353_));
 sky130_fd_sc_hd__mux2_1 _17124_ (.A0(\core.cpuregs[30][5] ),
    .A1(\core.cpuregs[31][5] ),
    .S(_10353_),
    .X(_10354_));
 sky130_fd_sc_hd__clkbuf_2 _17125_ (.A(_04649_),
    .X(_10355_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(_10351_),
    .A1(_10354_),
    .S(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__clkbuf_4 _17127_ (.A(_04539_),
    .X(_10357_));
 sky130_fd_sc_hd__clkbuf_2 _17128_ (.A(_10357_),
    .X(_10358_));
 sky130_fd_sc_hd__nand2_1 _17129_ (.A(_10356_),
    .B(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__clkbuf_2 _17130_ (.A(_10338_),
    .X(_10360_));
 sky130_fd_sc_hd__mux2_1 _17131_ (.A0(\core.cpuregs[12][5] ),
    .A1(\core.cpuregs[13][5] ),
    .S(_10360_),
    .X(_10361_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17132_ (.A(_04520_),
    .X(_10362_));
 sky130_fd_sc_hd__clkbuf_2 _17133_ (.A(_10362_),
    .X(_10363_));
 sky130_fd_sc_hd__mux2_1 _17134_ (.A0(\core.cpuregs[14][5] ),
    .A1(\core.cpuregs[15][5] ),
    .S(_10363_),
    .X(_10364_));
 sky130_fd_sc_hd__clkbuf_2 _17135_ (.A(_04528_),
    .X(_10365_));
 sky130_fd_sc_hd__clkbuf_2 _17136_ (.A(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__mux2_1 _17137_ (.A0(_10361_),
    .A1(_10364_),
    .S(_10366_),
    .X(_10367_));
 sky130_fd_sc_hd__clkbuf_8 _17138_ (.A(_04570_),
    .X(_10368_));
 sky130_fd_sc_hd__buf_1 _17139_ (.A(_10368_),
    .X(_10369_));
 sky130_fd_sc_hd__nand2_1 _17140_ (.A(_10367_),
    .B(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__clkbuf_2 _17141_ (.A(_04520_),
    .X(_10371_));
 sky130_fd_sc_hd__buf_2 _17142_ (.A(_10371_),
    .X(_10372_));
 sky130_fd_sc_hd__mux2_1 _17143_ (.A0(\core.cpuregs[8][5] ),
    .A1(\core.cpuregs[9][5] ),
    .S(_10372_),
    .X(_10373_));
 sky130_fd_sc_hd__clkbuf_2 _17144_ (.A(_04521_),
    .X(_10374_));
 sky130_fd_sc_hd__mux2_1 _17145_ (.A0(\core.cpuregs[10][5] ),
    .A1(\core.cpuregs[11][5] ),
    .S(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__clkbuf_2 _17146_ (.A(_10365_),
    .X(_10376_));
 sky130_fd_sc_hd__mux2_1 _17147_ (.A0(_10373_),
    .A1(_10375_),
    .S(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_10377_),
    .B(_10347_),
    .Y(_10378_));
 sky130_fd_sc_hd__inv_2 _17149_ (.A(_00004_),
    .Y(_10379_));
 sky130_fd_sc_hd__clkbuf_4 _17150_ (.A(_10379_),
    .X(_10380_));
 sky130_fd_sc_hd__and3_1 _17151_ (.A(_10370_),
    .B(_10378_),
    .C(_10380_),
    .X(_10381_));
 sky130_fd_sc_hd__a31o_1 _17152_ (.A1(_10337_),
    .A2(_10349_),
    .A3(_10359_),
    .B1(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__clkbuf_2 _17153_ (.A(_04552_),
    .X(_10383_));
 sky130_fd_sc_hd__buf_2 _17154_ (.A(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__nand2_2 _17155_ (.A(_04582_),
    .B(_04473_),
    .Y(_10385_));
 sky130_fd_sc_hd__clkbuf_2 _17156_ (.A(_10385_),
    .X(_10386_));
 sky130_fd_sc_hd__buf_2 _17157_ (.A(_10386_),
    .X(_10387_));
 sky130_fd_sc_hd__a21oi_2 _17158_ (.A1(_10382_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17159_ (.A(_10336_),
    .X(_10389_));
 sky130_fd_sc_hd__clkbuf_2 _17160_ (.A(_10339_),
    .X(_10390_));
 sky130_fd_sc_hd__mux2_1 _17161_ (.A0(\core.cpuregs[16][5] ),
    .A1(\core.cpuregs[17][5] ),
    .S(_10390_),
    .X(_10391_));
 sky130_fd_sc_hd__clkbuf_2 _17162_ (.A(_10371_),
    .X(_10392_));
 sky130_fd_sc_hd__buf_4 _17163_ (.A(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__mux2_1 _17164_ (.A0(\core.cpuregs[18][5] ),
    .A1(\core.cpuregs[19][5] ),
    .S(_10393_),
    .X(_10394_));
 sky130_fd_sc_hd__clkbuf_2 _17165_ (.A(_04640_),
    .X(_10395_));
 sky130_fd_sc_hd__clkbuf_2 _17166_ (.A(_10395_),
    .X(_10396_));
 sky130_fd_sc_hd__mux2_1 _17167_ (.A0(_10391_),
    .A1(_10394_),
    .S(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__buf_1 _17168_ (.A(_04549_),
    .X(_10398_));
 sky130_fd_sc_hd__buf_1 _17169_ (.A(_10398_),
    .X(_10399_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17170_ (.A(_10399_),
    .X(_10400_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(_10397_),
    .B(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__clkbuf_2 _17172_ (.A(_10392_),
    .X(_10402_));
 sky130_fd_sc_hd__mux2_1 _17173_ (.A0(\core.cpuregs[22][5] ),
    .A1(\core.cpuregs[23][5] ),
    .S(_10402_),
    .X(_10403_));
 sky130_fd_sc_hd__clkbuf_2 _17174_ (.A(_04522_),
    .X(_10404_));
 sky130_fd_sc_hd__mux2_1 _17175_ (.A0(\core.cpuregs[20][5] ),
    .A1(\core.cpuregs[21][5] ),
    .S(_10404_),
    .X(_10405_));
 sky130_fd_sc_hd__clkbuf_2 _17176_ (.A(_04537_),
    .X(_10406_));
 sky130_fd_sc_hd__mux2_2 _17177_ (.A0(_10403_),
    .A1(_10405_),
    .S(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17178_ (.A(_10369_),
    .X(_10408_));
 sky130_fd_sc_hd__nand2_1 _17179_ (.A(_10407_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__clkbuf_2 _17180_ (.A(_10357_),
    .X(_10410_));
 sky130_fd_sc_hd__clkbuf_2 _17181_ (.A(_10352_),
    .X(_10411_));
 sky130_fd_sc_hd__mux2_1 _17182_ (.A0(\core.cpuregs[6][5] ),
    .A1(\core.cpuregs[7][5] ),
    .S(_10411_),
    .X(_10412_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17183_ (.A(_04531_),
    .X(_10413_));
 sky130_fd_sc_hd__clkbuf_2 _17184_ (.A(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__mux2_1 _17185_ (.A0(\core.cpuregs[4][5] ),
    .A1(\core.cpuregs[5][5] ),
    .S(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__buf_4 _17186_ (.A(_04560_),
    .X(_10416_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(_10412_),
    .A1(_10415_),
    .S(_10416_),
    .X(_10417_));
 sky130_fd_sc_hd__buf_1 _17188_ (.A(_00004_),
    .X(_10418_));
 sky130_fd_sc_hd__clkbuf_2 _17189_ (.A(_10418_),
    .X(_10419_));
 sky130_fd_sc_hd__clkbuf_2 _17190_ (.A(_09613_),
    .X(_10420_));
 sky130_fd_sc_hd__mux2_1 _17191_ (.A0(\core.cpuregs[0][5] ),
    .A1(\core.cpuregs[1][5] ),
    .S(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__clkbuf_2 _17192_ (.A(_10338_),
    .X(_10422_));
 sky130_fd_sc_hd__mux2_1 _17193_ (.A0(\core.cpuregs[2][5] ),
    .A1(\core.cpuregs[3][5] ),
    .S(_10422_),
    .X(_10423_));
 sky130_fd_sc_hd__clkbuf_2 _17194_ (.A(_09650_),
    .X(_10424_));
 sky130_fd_sc_hd__mux2_2 _17195_ (.A0(_10421_),
    .A1(_10423_),
    .S(_10424_),
    .X(_10425_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17196_ (.A(_10398_),
    .X(_10426_));
 sky130_fd_sc_hd__and2_1 _17197_ (.A(_10425_),
    .B(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__a211oi_2 _17198_ (.A1(_10410_),
    .A2(_10417_),
    .B1(_10419_),
    .C1(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__a31o_1 _17199_ (.A1(_10389_),
    .A2(_10401_),
    .A3(_10409_),
    .B1(_10428_),
    .X(_10429_));
 sky130_fd_sc_hd__inv_2 _17200_ (.A(_04656_),
    .Y(_10430_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17201_ (.A(_10430_),
    .X(_10431_));
 sky130_fd_sc_hd__nand2_1 _17202_ (.A(_10429_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__a22o_1 _17203_ (.A1(\core.decoded_imm[5] ),
    .A2(_10318_),
    .B1(_10388_),
    .B2(_10432_),
    .X(_10433_));
 sky130_fd_sc_hd__clkbuf_4 _17204_ (.A(_10321_),
    .X(_10434_));
 sky130_fd_sc_hd__mux2_1 _17205_ (.A0(_10433_),
    .A1(_04714_),
    .S(_10434_),
    .X(_10435_));
 sky130_fd_sc_hd__clkbuf_2 _17206_ (.A(_10435_),
    .X(_00609_));
 sky130_fd_sc_hd__clkbuf_4 _17207_ (.A(_04496_),
    .X(_10436_));
 sky130_fd_sc_hd__mux2_2 _17208_ (.A0(\core.cpuregs[24][6] ),
    .A1(\core.cpuregs[25][6] ),
    .S(_10340_),
    .X(_10437_));
 sky130_fd_sc_hd__mux2_1 _17209_ (.A0(\core.cpuregs[26][6] ),
    .A1(\core.cpuregs[27][6] ),
    .S(_10342_),
    .X(_10438_));
 sky130_fd_sc_hd__mux2_1 _17210_ (.A0(_10437_),
    .A1(_10438_),
    .S(_10344_),
    .X(_10439_));
 sky130_fd_sc_hd__nand2_1 _17211_ (.A(_10439_),
    .B(_10348_),
    .Y(_10440_));
 sky130_fd_sc_hd__mux2_1 _17212_ (.A0(\core.cpuregs[28][6] ),
    .A1(\core.cpuregs[29][6] ),
    .S(_10350_),
    .X(_10441_));
 sky130_fd_sc_hd__mux2_1 _17213_ (.A0(\core.cpuregs[30][6] ),
    .A1(\core.cpuregs[31][6] ),
    .S(_10353_),
    .X(_10442_));
 sky130_fd_sc_hd__mux2_1 _17214_ (.A0(_10441_),
    .A1(_10442_),
    .S(_10355_),
    .X(_10443_));
 sky130_fd_sc_hd__nand2_2 _17215_ (.A(_10443_),
    .B(_10358_),
    .Y(_10444_));
 sky130_fd_sc_hd__mux2_1 _17216_ (.A0(\core.cpuregs[12][6] ),
    .A1(\core.cpuregs[13][6] ),
    .S(_10360_),
    .X(_10445_));
 sky130_fd_sc_hd__buf_2 _17217_ (.A(_10362_),
    .X(_10446_));
 sky130_fd_sc_hd__mux2_1 _17218_ (.A0(\core.cpuregs[14][6] ),
    .A1(\core.cpuregs[15][6] ),
    .S(_10446_),
    .X(_10447_));
 sky130_fd_sc_hd__mux2_1 _17219_ (.A0(_10445_),
    .A1(_10447_),
    .S(_10366_),
    .X(_10448_));
 sky130_fd_sc_hd__clkbuf_8 _17220_ (.A(_10368_),
    .X(_10449_));
 sky130_fd_sc_hd__nand2_1 _17221_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__mux2_1 _17222_ (.A0(\core.cpuregs[8][6] ),
    .A1(\core.cpuregs[9][6] ),
    .S(_10372_),
    .X(_10451_));
 sky130_fd_sc_hd__mux2_1 _17223_ (.A0(\core.cpuregs[10][6] ),
    .A1(\core.cpuregs[11][6] ),
    .S(_10374_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _17224_ (.A0(_10451_),
    .A1(_01575_),
    .S(_10376_),
    .X(_01576_));
 sky130_fd_sc_hd__nand2_1 _17225_ (.A(_01576_),
    .B(_10347_),
    .Y(_01577_));
 sky130_fd_sc_hd__and3_1 _17226_ (.A(_10450_),
    .B(_01577_),
    .C(_10380_),
    .X(_01578_));
 sky130_fd_sc_hd__a31o_1 _17227_ (.A1(_10337_),
    .A2(_10440_),
    .A3(_10444_),
    .B1(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__a21oi_4 _17228_ (.A1(_01579_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_01580_));
 sky130_fd_sc_hd__mux2_1 _17229_ (.A0(\core.cpuregs[16][6] ),
    .A1(\core.cpuregs[17][6] ),
    .S(_10390_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _17230_ (.A0(\core.cpuregs[18][6] ),
    .A1(\core.cpuregs[19][6] ),
    .S(_10393_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _17231_ (.A0(_01581_),
    .A1(_01582_),
    .S(_10396_),
    .X(_01583_));
 sky130_fd_sc_hd__nand2_1 _17232_ (.A(_01583_),
    .B(_10400_),
    .Y(_01584_));
 sky130_fd_sc_hd__mux2_1 _17233_ (.A0(\core.cpuregs[22][6] ),
    .A1(\core.cpuregs[23][6] ),
    .S(_10402_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _17234_ (.A0(\core.cpuregs[20][6] ),
    .A1(\core.cpuregs[21][6] ),
    .S(_10404_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _17235_ (.A0(_01585_),
    .A1(_01586_),
    .S(_10406_),
    .X(_01587_));
 sky130_fd_sc_hd__nand2_1 _17236_ (.A(_01587_),
    .B(_10408_),
    .Y(_01588_));
 sky130_fd_sc_hd__mux2_1 _17237_ (.A0(\core.cpuregs[6][6] ),
    .A1(\core.cpuregs[7][6] ),
    .S(_10411_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _17238_ (.A0(\core.cpuregs[4][6] ),
    .A1(\core.cpuregs[5][6] ),
    .S(_10414_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _17239_ (.A0(_01589_),
    .A1(_01590_),
    .S(_10416_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _17240_ (.A0(\core.cpuregs[0][6] ),
    .A1(\core.cpuregs[1][6] ),
    .S(_10420_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(\core.cpuregs[2][6] ),
    .A1(\core.cpuregs[3][6] ),
    .S(_10422_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _17242_ (.A0(_01592_),
    .A1(_01593_),
    .S(_10424_),
    .X(_01594_));
 sky130_fd_sc_hd__and2_1 _17243_ (.A(_01594_),
    .B(_10426_),
    .X(_01595_));
 sky130_fd_sc_hd__a211oi_1 _17244_ (.A1(_10410_),
    .A2(_01591_),
    .B1(_10419_),
    .C1(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__a31o_2 _17245_ (.A1(_10389_),
    .A2(_01584_),
    .A3(_01588_),
    .B1(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__nand2_1 _17246_ (.A(_01597_),
    .B(_10431_),
    .Y(_01598_));
 sky130_fd_sc_hd__a22o_1 _17247_ (.A1(\core.decoded_imm[6] ),
    .A2(_10436_),
    .B1(_01580_),
    .B2(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _17248_ (.A0(_01599_),
    .A1(_04709_),
    .S(_10434_),
    .X(_01600_));
 sky130_fd_sc_hd__clkbuf_1 _17249_ (.A(_01600_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _17250_ (.A0(\core.cpuregs[24][7] ),
    .A1(\core.cpuregs[25][7] ),
    .S(_10340_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _17251_ (.A0(\core.cpuregs[26][7] ),
    .A1(\core.cpuregs[27][7] ),
    .S(_10342_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _17252_ (.A0(_01601_),
    .A1(_01602_),
    .S(_10344_),
    .X(_01603_));
 sky130_fd_sc_hd__nand2_1 _17253_ (.A(_01603_),
    .B(_10348_),
    .Y(_01604_));
 sky130_fd_sc_hd__mux2_1 _17254_ (.A0(\core.cpuregs[28][7] ),
    .A1(\core.cpuregs[29][7] ),
    .S(_10350_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _17255_ (.A0(\core.cpuregs[30][7] ),
    .A1(\core.cpuregs[31][7] ),
    .S(_10353_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _17256_ (.A0(_01605_),
    .A1(_01606_),
    .S(_10355_),
    .X(_01607_));
 sky130_fd_sc_hd__buf_2 _17257_ (.A(_10357_),
    .X(_01608_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(_01607_),
    .B(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__buf_2 _17259_ (.A(_10362_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _17260_ (.A0(\core.cpuregs[12][7] ),
    .A1(\core.cpuregs[13][7] ),
    .S(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _17261_ (.A0(\core.cpuregs[14][7] ),
    .A1(\core.cpuregs[15][7] ),
    .S(_10446_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_2 _17262_ (.A0(_01611_),
    .A1(_01612_),
    .S(_10366_),
    .X(_01613_));
 sky130_fd_sc_hd__nand2_4 _17263_ (.A(_01613_),
    .B(_10449_),
    .Y(_01614_));
 sky130_fd_sc_hd__mux2_1 _17264_ (.A0(\core.cpuregs[8][7] ),
    .A1(\core.cpuregs[9][7] ),
    .S(_10372_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _17265_ (.A0(\core.cpuregs[10][7] ),
    .A1(\core.cpuregs[11][7] ),
    .S(_10374_),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_2 _17266_ (.A0(_01615_),
    .A1(_01616_),
    .S(_10376_),
    .X(_01617_));
 sky130_fd_sc_hd__clkbuf_4 _17267_ (.A(_10346_),
    .X(_01618_));
 sky130_fd_sc_hd__nand2_4 _17268_ (.A(_01617_),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__and3_1 _17269_ (.A(_01614_),
    .B(_01619_),
    .C(_10380_),
    .X(_01620_));
 sky130_fd_sc_hd__a31o_1 _17270_ (.A1(_10337_),
    .A2(_01604_),
    .A3(_01609_),
    .B1(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__a21oi_2 _17271_ (.A1(_01621_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_01622_));
 sky130_fd_sc_hd__mux2_1 _17272_ (.A0(\core.cpuregs[16][7] ),
    .A1(\core.cpuregs[17][7] ),
    .S(_10390_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_2 _17273_ (.A0(\core.cpuregs[18][7] ),
    .A1(\core.cpuregs[19][7] ),
    .S(_10393_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _17274_ (.A0(_01623_),
    .A1(_01624_),
    .S(_10396_),
    .X(_01625_));
 sky130_fd_sc_hd__nand2_1 _17275_ (.A(_01625_),
    .B(_10400_),
    .Y(_01626_));
 sky130_fd_sc_hd__mux2_1 _17276_ (.A0(\core.cpuregs[22][7] ),
    .A1(\core.cpuregs[23][7] ),
    .S(_10402_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _17277_ (.A0(\core.cpuregs[20][7] ),
    .A1(\core.cpuregs[21][7] ),
    .S(_10404_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _17278_ (.A0(_01627_),
    .A1(_01628_),
    .S(_10406_),
    .X(_01629_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17279_ (.A(_10369_),
    .X(_01630_));
 sky130_fd_sc_hd__nand2_1 _17280_ (.A(_01629_),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__clkbuf_2 _17281_ (.A(_04539_),
    .X(_01632_));
 sky130_fd_sc_hd__clkbuf_2 _17282_ (.A(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _17283_ (.A0(\core.cpuregs[6][7] ),
    .A1(\core.cpuregs[7][7] ),
    .S(_10411_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _17284_ (.A0(\core.cpuregs[4][7] ),
    .A1(\core.cpuregs[5][7] ),
    .S(_10414_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _17285_ (.A0(_01634_),
    .A1(_01635_),
    .S(_10416_),
    .X(_01636_));
 sky130_fd_sc_hd__clkbuf_2 _17286_ (.A(_09648_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _17287_ (.A0(\core.cpuregs[0][7] ),
    .A1(\core.cpuregs[1][7] ),
    .S(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__clkbuf_2 _17288_ (.A(_10338_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _17289_ (.A0(\core.cpuregs[2][7] ),
    .A1(\core.cpuregs[3][7] ),
    .S(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _17290_ (.A0(_01638_),
    .A1(_01640_),
    .S(_10424_),
    .X(_01641_));
 sky130_fd_sc_hd__buf_1 _17291_ (.A(_10346_),
    .X(_01642_));
 sky130_fd_sc_hd__and2_1 _17292_ (.A(_01641_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__a211oi_1 _17293_ (.A1(_01633_),
    .A2(_01636_),
    .B1(_10419_),
    .C1(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__a31o_1 _17294_ (.A1(_10389_),
    .A2(_01626_),
    .A3(_01631_),
    .B1(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__nand2_1 _17295_ (.A(_01645_),
    .B(_10431_),
    .Y(_01646_));
 sky130_fd_sc_hd__a22o_1 _17296_ (.A1(\core.decoded_imm[7] ),
    .A2(_10436_),
    .B1(_01622_),
    .B2(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _17297_ (.A0(_01647_),
    .A1(_04705_),
    .S(_10434_),
    .X(_01648_));
 sky130_fd_sc_hd__clkbuf_1 _17298_ (.A(_01648_),
    .X(_00611_));
 sky130_fd_sc_hd__inv_2 _17299_ (.A(_10322_),
    .Y(_01649_));
 sky130_fd_sc_hd__o21ai_1 _17300_ (.A1(_06131_),
    .A2(_04474_),
    .B1(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__clkbuf_4 _17301_ (.A(_10389_),
    .X(_01651_));
 sky130_fd_sc_hd__clkbuf_4 _17302_ (.A(_10340_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _17303_ (.A0(\core.cpuregs[16][8] ),
    .A1(\core.cpuregs[17][8] ),
    .S(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_4 _17304_ (.A0(\core.cpuregs[18][8] ),
    .A1(\core.cpuregs[19][8] ),
    .S(_01652_),
    .X(_01654_));
 sky130_fd_sc_hd__clkbuf_2 _17305_ (.A(_10424_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _17306_ (.A0(_01653_),
    .A1(_01654_),
    .S(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17307_ (.A(_10348_),
    .X(_01657_));
 sky130_fd_sc_hd__nand2_1 _17308_ (.A(_01656_),
    .B(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__buf_4 _17309_ (.A(_10340_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _17310_ (.A0(\core.cpuregs[22][8] ),
    .A1(\core.cpuregs[23][8] ),
    .S(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_4 _17311_ (.A0(\core.cpuregs[20][8] ),
    .A1(\core.cpuregs[21][8] ),
    .S(_01659_),
    .X(_01661_));
 sky130_fd_sc_hd__clkbuf_2 _17312_ (.A(_04537_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _17313_ (.A0(_01660_),
    .A1(_01661_),
    .S(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17314_ (.A(_10408_),
    .X(_01664_));
 sky130_fd_sc_hd__nand2_1 _17315_ (.A(_01663_),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__clkbuf_2 _17316_ (.A(_10420_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(\core.cpuregs[6][8] ),
    .A1(\core.cpuregs[7][8] ),
    .S(_01666_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_2 _17318_ (.A0(\core.cpuregs[4][8] ),
    .A1(\core.cpuregs[5][8] ),
    .S(_01666_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _17319_ (.A0(_01667_),
    .A1(_01668_),
    .S(_01662_),
    .X(_01669_));
 sky130_fd_sc_hd__clkbuf_4 _17320_ (.A(_10371_),
    .X(_01670_));
 sky130_fd_sc_hd__clkbuf_2 _17321_ (.A(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _17322_ (.A0(\core.cpuregs[0][8] ),
    .A1(\core.cpuregs[1][8] ),
    .S(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(\core.cpuregs[2][8] ),
    .A1(\core.cpuregs[3][8] ),
    .S(_01671_),
    .X(_01673_));
 sky130_fd_sc_hd__clkbuf_2 _17324_ (.A(_10376_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _17325_ (.A0(_01672_),
    .A1(_01673_),
    .S(_01674_),
    .X(_01675_));
 sky130_fd_sc_hd__clkbuf_4 _17326_ (.A(_10399_),
    .X(_01676_));
 sky130_fd_sc_hd__and2_1 _17327_ (.A(_01675_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__a211oi_1 _17328_ (.A1(_01664_),
    .A2(_01669_),
    .B1(_01651_),
    .C1(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__a31o_1 _17329_ (.A1(_01651_),
    .A2(_01658_),
    .A3(_01665_),
    .B1(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__clkbuf_4 _17330_ (.A(_10336_),
    .X(_01680_));
 sky130_fd_sc_hd__clkbuf_2 _17331_ (.A(_10420_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _17332_ (.A0(\core.cpuregs[24][8] ),
    .A1(\core.cpuregs[25][8] ),
    .S(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _17333_ (.A0(\core.cpuregs[26][8] ),
    .A1(\core.cpuregs[27][8] ),
    .S(_01681_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _17334_ (.A0(_01682_),
    .A1(_01683_),
    .S(_01655_),
    .X(_01684_));
 sky130_fd_sc_hd__nand2_1 _17335_ (.A(_01684_),
    .B(_01657_),
    .Y(_01685_));
 sky130_fd_sc_hd__clkbuf_4 _17336_ (.A(_10363_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _17337_ (.A0(\core.cpuregs[28][8] ),
    .A1(\core.cpuregs[29][8] ),
    .S(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _17338_ (.A0(\core.cpuregs[30][8] ),
    .A1(\core.cpuregs[31][8] ),
    .S(_01686_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _17339_ (.A0(_01687_),
    .A1(_01688_),
    .S(_01674_),
    .X(_01689_));
 sky130_fd_sc_hd__nand2_1 _17340_ (.A(_01689_),
    .B(_10408_),
    .Y(_01690_));
 sky130_fd_sc_hd__clkbuf_2 _17341_ (.A(_10339_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _17342_ (.A0(\core.cpuregs[8][8] ),
    .A1(\core.cpuregs[9][8] ),
    .S(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\core.cpuregs[10][8] ),
    .A1(\core.cpuregs[11][8] ),
    .S(_01691_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _17344_ (.A0(_01692_),
    .A1(_01693_),
    .S(_10396_),
    .X(_01694_));
 sky130_fd_sc_hd__clkbuf_2 _17345_ (.A(_04638_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _17346_ (.A0(\core.cpuregs[12][8] ),
    .A1(\core.cpuregs[13][8] ),
    .S(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(\core.cpuregs[14][8] ),
    .A1(\core.cpuregs[15][8] ),
    .S(_01695_),
    .X(_01697_));
 sky130_fd_sc_hd__clkbuf_2 _17348_ (.A(_04641_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _17349_ (.A0(_01696_),
    .A1(_01697_),
    .S(_01698_),
    .X(_01699_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17350_ (.A(_10368_),
    .X(_01700_));
 sky130_fd_sc_hd__and2_2 _17351_ (.A(_01699_),
    .B(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__a211oi_2 _17352_ (.A1(_01676_),
    .A2(_01694_),
    .B1(_01680_),
    .C1(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__a31o_1 _17353_ (.A1(_01680_),
    .A2(_01685_),
    .A3(_01690_),
    .B1(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__a21oi_1 _17354_ (.A1(_01703_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_01704_));
 sky130_fd_sc_hd__a21boi_1 _17355_ (.A1(_10431_),
    .A2(_01679_),
    .B1_N(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__o22a_1 _17356_ (.A1(\core.pcpi_rs2[8] ),
    .A2(_01649_),
    .B1(_01650_),
    .B2(_01705_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _17357_ (.A0(\core.cpuregs[24][9] ),
    .A1(\core.cpuregs[25][9] ),
    .S(_10340_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _17358_ (.A0(\core.cpuregs[26][9] ),
    .A1(\core.cpuregs[27][9] ),
    .S(_10342_),
    .X(_01707_));
 sky130_fd_sc_hd__clkbuf_2 _17359_ (.A(_04641_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _17360_ (.A0(_01706_),
    .A1(_01707_),
    .S(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__nand2_2 _17361_ (.A(_01709_),
    .B(_10348_),
    .Y(_01710_));
 sky130_fd_sc_hd__mux2_1 _17362_ (.A0(\core.cpuregs[28][9] ),
    .A1(\core.cpuregs[29][9] ),
    .S(_10350_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _17363_ (.A0(\core.cpuregs[30][9] ),
    .A1(\core.cpuregs[31][9] ),
    .S(_10353_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _17364_ (.A0(_01711_),
    .A1(_01712_),
    .S(_10355_),
    .X(_01713_));
 sky130_fd_sc_hd__nand2_2 _17365_ (.A(_01713_),
    .B(_01608_),
    .Y(_01714_));
 sky130_fd_sc_hd__mux2_1 _17366_ (.A0(\core.cpuregs[12][9] ),
    .A1(\core.cpuregs[13][9] ),
    .S(_01610_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _17367_ (.A0(\core.cpuregs[14][9] ),
    .A1(\core.cpuregs[15][9] ),
    .S(_10446_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_2 _17368_ (.A0(_01715_),
    .A1(_01716_),
    .S(_10366_),
    .X(_01717_));
 sky130_fd_sc_hd__nand2_4 _17369_ (.A(_01717_),
    .B(_10449_),
    .Y(_01718_));
 sky130_fd_sc_hd__mux2_1 _17370_ (.A0(\core.cpuregs[8][9] ),
    .A1(\core.cpuregs[9][9] ),
    .S(_10372_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _17371_ (.A0(\core.cpuregs[10][9] ),
    .A1(\core.cpuregs[11][9] ),
    .S(_10374_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _17372_ (.A0(_01719_),
    .A1(_01720_),
    .S(_10376_),
    .X(_01721_));
 sky130_fd_sc_hd__nand2_1 _17373_ (.A(_01721_),
    .B(_01618_),
    .Y(_01722_));
 sky130_fd_sc_hd__and3_1 _17374_ (.A(_01718_),
    .B(_01722_),
    .C(_10380_),
    .X(_01723_));
 sky130_fd_sc_hd__a31o_1 _17375_ (.A1(_10337_),
    .A2(_01710_),
    .A3(_01714_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__buf_4 _17376_ (.A(_10383_),
    .X(_01725_));
 sky130_fd_sc_hd__buf_4 _17377_ (.A(_10386_),
    .X(_01726_));
 sky130_fd_sc_hd__a21oi_2 _17378_ (.A1(_01724_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__mux2_1 _17379_ (.A0(\core.cpuregs[16][9] ),
    .A1(\core.cpuregs[17][9] ),
    .S(_10390_),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _17380_ (.A0(\core.cpuregs[18][9] ),
    .A1(\core.cpuregs[19][9] ),
    .S(_10393_),
    .X(_01729_));
 sky130_fd_sc_hd__clkbuf_2 _17381_ (.A(_10395_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _17382_ (.A0(_01728_),
    .A1(_01729_),
    .S(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_2 _17383_ (.A(_01731_),
    .B(_10400_),
    .Y(_01732_));
 sky130_fd_sc_hd__mux2_1 _17384_ (.A0(\core.cpuregs[22][9] ),
    .A1(\core.cpuregs[23][9] ),
    .S(_10402_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _17385_ (.A0(\core.cpuregs[20][9] ),
    .A1(\core.cpuregs[21][9] ),
    .S(_10404_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_2 _17386_ (.A0(_01733_),
    .A1(_01734_),
    .S(_10406_),
    .X(_01735_));
 sky130_fd_sc_hd__nand2_1 _17387_ (.A(_01735_),
    .B(_01630_),
    .Y(_01736_));
 sky130_fd_sc_hd__mux2_1 _17388_ (.A0(\core.cpuregs[6][9] ),
    .A1(\core.cpuregs[7][9] ),
    .S(_10411_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_2 _17389_ (.A0(\core.cpuregs[4][9] ),
    .A1(\core.cpuregs[5][9] ),
    .S(_10414_),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _17390_ (.A0(_01737_),
    .A1(_01738_),
    .S(_10416_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _17391_ (.A0(\core.cpuregs[0][9] ),
    .A1(\core.cpuregs[1][9] ),
    .S(_01637_),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _17392_ (.A0(\core.cpuregs[2][9] ),
    .A1(\core.cpuregs[3][9] ),
    .S(_01639_),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _17393_ (.A0(_01740_),
    .A1(_01741_),
    .S(_10424_),
    .X(_01742_));
 sky130_fd_sc_hd__and2_1 _17394_ (.A(_01742_),
    .B(_01642_),
    .X(_01743_));
 sky130_fd_sc_hd__a211oi_2 _17395_ (.A1(_01633_),
    .A2(_01739_),
    .B1(_10419_),
    .C1(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a31o_1 _17396_ (.A1(_10389_),
    .A2(_01732_),
    .A3(_01736_),
    .B1(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__buf_2 _17397_ (.A(_10430_),
    .X(_01746_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17398_ (.A(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(_01745_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__a22o_1 _17400_ (.A1(\core.decoded_imm[9] ),
    .A2(_10436_),
    .B1(_01727_),
    .B2(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_4 _17401_ (.A0(_01749_),
    .A1(\core.pcpi_rs2[9] ),
    .S(_10434_),
    .X(_01750_));
 sky130_fd_sc_hd__clkbuf_1 _17402_ (.A(_01750_),
    .X(_00613_));
 sky130_fd_sc_hd__clkbuf_2 _17403_ (.A(_04567_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _17404_ (.A0(\core.cpuregs[24][10] ),
    .A1(\core.cpuregs[25][10] ),
    .S(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__clkbuf_2 _17405_ (.A(_04636_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _17406_ (.A0(\core.cpuregs[26][10] ),
    .A1(\core.cpuregs[27][10] ),
    .S(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _17407_ (.A0(_01752_),
    .A1(_01754_),
    .S(_01708_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_01755_),
    .B(_10348_),
    .Y(_01756_));
 sky130_fd_sc_hd__buf_4 _17409_ (.A(_04662_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _17410_ (.A0(\core.cpuregs[28][10] ),
    .A1(\core.cpuregs[29][10] ),
    .S(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__clkbuf_2 _17411_ (.A(_10352_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _17412_ (.A0(\core.cpuregs[30][10] ),
    .A1(\core.cpuregs[31][10] ),
    .S(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _17413_ (.A0(_01758_),
    .A1(_01760_),
    .S(_10355_),
    .X(_01761_));
 sky130_fd_sc_hd__nand2_1 _17414_ (.A(_01761_),
    .B(_01608_),
    .Y(_01762_));
 sky130_fd_sc_hd__mux2_1 _17415_ (.A0(\core.cpuregs[12][10] ),
    .A1(\core.cpuregs[13][10] ),
    .S(_01610_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _17416_ (.A0(\core.cpuregs[14][10] ),
    .A1(\core.cpuregs[15][10] ),
    .S(_10446_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _17417_ (.A0(_01763_),
    .A1(_01764_),
    .S(_10366_),
    .X(_01765_));
 sky130_fd_sc_hd__nand2_1 _17418_ (.A(_01765_),
    .B(_10449_),
    .Y(_01766_));
 sky130_fd_sc_hd__mux2_1 _17419_ (.A0(\core.cpuregs[8][10] ),
    .A1(\core.cpuregs[9][10] ),
    .S(_10372_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _17420_ (.A0(\core.cpuregs[10][10] ),
    .A1(\core.cpuregs[11][10] ),
    .S(_10374_),
    .X(_01768_));
 sky130_fd_sc_hd__clkbuf_2 _17421_ (.A(_04640_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _17422_ (.A0(_01767_),
    .A1(_01768_),
    .S(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_2 _17423_ (.A(_01770_),
    .B(_01618_),
    .Y(_01771_));
 sky130_fd_sc_hd__and3_1 _17424_ (.A(_01766_),
    .B(_01771_),
    .C(_10380_),
    .X(_01772_));
 sky130_fd_sc_hd__a31o_1 _17425_ (.A1(_10337_),
    .A2(_01756_),
    .A3(_01762_),
    .B1(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__a21oi_2 _17426_ (.A1(_01773_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01774_));
 sky130_fd_sc_hd__mux2_1 _17427_ (.A0(\core.cpuregs[16][10] ),
    .A1(\core.cpuregs[17][10] ),
    .S(_10390_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _17428_ (.A0(\core.cpuregs[18][10] ),
    .A1(\core.cpuregs[19][10] ),
    .S(_10393_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _17429_ (.A0(_01775_),
    .A1(_01776_),
    .S(_01730_),
    .X(_01777_));
 sky130_fd_sc_hd__nand2_1 _17430_ (.A(_01777_),
    .B(_10400_),
    .Y(_01778_));
 sky130_fd_sc_hd__mux2_2 _17431_ (.A0(\core.cpuregs[22][10] ),
    .A1(\core.cpuregs[23][10] ),
    .S(_10402_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _17432_ (.A0(\core.cpuregs[20][10] ),
    .A1(\core.cpuregs[21][10] ),
    .S(_10404_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(_01779_),
    .A1(_01780_),
    .S(_10406_),
    .X(_01781_));
 sky130_fd_sc_hd__nand2_1 _17434_ (.A(_01781_),
    .B(_01630_),
    .Y(_01782_));
 sky130_fd_sc_hd__clkbuf_2 _17435_ (.A(_10352_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _17436_ (.A0(\core.cpuregs[6][10] ),
    .A1(\core.cpuregs[7][10] ),
    .S(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__clkbuf_2 _17437_ (.A(_10413_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _17438_ (.A0(\core.cpuregs[4][10] ),
    .A1(\core.cpuregs[5][10] ),
    .S(_01785_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _17439_ (.A0(_01784_),
    .A1(_01786_),
    .S(_10416_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_8 _17440_ (.A0(\core.cpuregs[0][10] ),
    .A1(\core.cpuregs[1][10] ),
    .S(_01637_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _17441_ (.A0(\core.cpuregs[2][10] ),
    .A1(\core.cpuregs[3][10] ),
    .S(_01639_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _17442_ (.A0(_01788_),
    .A1(_01789_),
    .S(_10424_),
    .X(_01790_));
 sky130_fd_sc_hd__and2_1 _17443_ (.A(_01790_),
    .B(_01642_),
    .X(_01791_));
 sky130_fd_sc_hd__a211oi_2 _17444_ (.A1(_01633_),
    .A2(_01787_),
    .B1(_10419_),
    .C1(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__a31o_1 _17445_ (.A1(_10389_),
    .A2(_01778_),
    .A3(_01782_),
    .B1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(_01793_),
    .B(_01747_),
    .Y(_01794_));
 sky130_fd_sc_hd__a22o_1 _17447_ (.A1(\core.decoded_imm[10] ),
    .A2(_10436_),
    .B1(_01774_),
    .B2(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _17448_ (.A0(_01795_),
    .A1(\core.pcpi_rs2[10] ),
    .S(_10434_),
    .X(_01796_));
 sky130_fd_sc_hd__clkbuf_2 _17449_ (.A(_01796_),
    .X(_00614_));
 sky130_fd_sc_hd__buf_2 _17450_ (.A(_10418_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _17451_ (.A0(\core.cpuregs[24][11] ),
    .A1(\core.cpuregs[25][11] ),
    .S(_01751_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _17452_ (.A0(\core.cpuregs[26][11] ),
    .A1(\core.cpuregs[27][11] ),
    .S(_01753_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _17453_ (.A0(_01798_),
    .A1(_01799_),
    .S(_01708_),
    .X(_01800_));
 sky130_fd_sc_hd__clkbuf_4 _17454_ (.A(_10347_),
    .X(_01801_));
 sky130_fd_sc_hd__nand2_1 _17455_ (.A(_01800_),
    .B(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__mux2_1 _17456_ (.A0(\core.cpuregs[28][11] ),
    .A1(\core.cpuregs[29][11] ),
    .S(_01757_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _17457_ (.A0(\core.cpuregs[30][11] ),
    .A1(\core.cpuregs[31][11] ),
    .S(_01759_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _17458_ (.A0(_01803_),
    .A1(_01804_),
    .S(_10355_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _17459_ (.A(_01805_),
    .B(_01608_),
    .Y(_01806_));
 sky130_fd_sc_hd__mux2_1 _17460_ (.A0(\core.cpuregs[12][11] ),
    .A1(\core.cpuregs[13][11] ),
    .S(_01610_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _17461_ (.A0(\core.cpuregs[14][11] ),
    .A1(\core.cpuregs[15][11] ),
    .S(_10446_),
    .X(_01808_));
 sky130_fd_sc_hd__buf_4 _17462_ (.A(_10365_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_2 _17463_ (.A0(_01807_),
    .A1(_01808_),
    .S(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__nand2_4 _17464_ (.A(_01810_),
    .B(_10449_),
    .Y(_01811_));
 sky130_fd_sc_hd__mux2_1 _17465_ (.A0(\core.cpuregs[8][11] ),
    .A1(\core.cpuregs[9][11] ),
    .S(_10372_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _17466_ (.A0(\core.cpuregs[10][11] ),
    .A1(\core.cpuregs[11][11] ),
    .S(_10374_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_2 _17467_ (.A0(_01812_),
    .A1(_01813_),
    .S(_01769_),
    .X(_01814_));
 sky130_fd_sc_hd__nand2_8 _17468_ (.A(_01814_),
    .B(_01618_),
    .Y(_01815_));
 sky130_fd_sc_hd__and3_1 _17469_ (.A(_01811_),
    .B(_01815_),
    .C(_10380_),
    .X(_01816_));
 sky130_fd_sc_hd__a31o_1 _17470_ (.A1(_01797_),
    .A2(_01802_),
    .A3(_01806_),
    .B1(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__a21oi_2 _17471_ (.A1(_01817_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01818_));
 sky130_fd_sc_hd__clkbuf_4 _17472_ (.A(_10336_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _17473_ (.A0(\core.cpuregs[16][11] ),
    .A1(\core.cpuregs[17][11] ),
    .S(_10390_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _17474_ (.A0(\core.cpuregs[18][11] ),
    .A1(\core.cpuregs[19][11] ),
    .S(_10393_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _17475_ (.A0(_01820_),
    .A1(_01821_),
    .S(_01730_),
    .X(_01822_));
 sky130_fd_sc_hd__nand2_1 _17476_ (.A(_01822_),
    .B(_10400_),
    .Y(_01823_));
 sky130_fd_sc_hd__mux2_1 _17477_ (.A0(\core.cpuregs[22][11] ),
    .A1(\core.cpuregs[23][11] ),
    .S(_10402_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _17478_ (.A0(\core.cpuregs[20][11] ),
    .A1(\core.cpuregs[21][11] ),
    .S(_10404_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _17479_ (.A0(_01824_),
    .A1(_01825_),
    .S(_10406_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _17480_ (.A(_01826_),
    .B(_01630_),
    .Y(_01827_));
 sky130_fd_sc_hd__mux2_1 _17481_ (.A0(\core.cpuregs[6][11] ),
    .A1(\core.cpuregs[7][11] ),
    .S(_01783_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_8 _17482_ (.A0(\core.cpuregs[4][11] ),
    .A1(\core.cpuregs[5][11] ),
    .S(_01785_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _17483_ (.A0(_01828_),
    .A1(_01829_),
    .S(_10416_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _17484_ (.A0(\core.cpuregs[0][11] ),
    .A1(\core.cpuregs[1][11] ),
    .S(_01637_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_8 _17485_ (.A0(\core.cpuregs[2][11] ),
    .A1(\core.cpuregs[3][11] ),
    .S(_01639_),
    .X(_01832_));
 sky130_fd_sc_hd__clkbuf_2 _17486_ (.A(_09650_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _17487_ (.A0(_01831_),
    .A1(_01832_),
    .S(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__and2_1 _17488_ (.A(_01834_),
    .B(_01642_),
    .X(_01835_));
 sky130_fd_sc_hd__a211oi_1 _17489_ (.A1(_01633_),
    .A2(_01830_),
    .B1(_10419_),
    .C1(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__a31o_1 _17490_ (.A1(_01819_),
    .A2(_01823_),
    .A3(_01827_),
    .B1(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__nand2_1 _17491_ (.A(_01837_),
    .B(_01747_),
    .Y(_01838_));
 sky130_fd_sc_hd__a22o_1 _17492_ (.A1(\core.decoded_imm[11] ),
    .A2(_10436_),
    .B1(_01818_),
    .B2(_01838_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_4 _17493_ (.A0(_01839_),
    .A1(\core.pcpi_rs2[11] ),
    .S(_10434_),
    .X(_01840_));
 sky130_fd_sc_hd__clkbuf_1 _17494_ (.A(_01840_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _17495_ (.A0(\core.cpuregs[24][12] ),
    .A1(\core.cpuregs[25][12] ),
    .S(_01751_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _17496_ (.A0(\core.cpuregs[26][12] ),
    .A1(\core.cpuregs[27][12] ),
    .S(_01753_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _17497_ (.A0(_01841_),
    .A1(_01842_),
    .S(_01708_),
    .X(_01843_));
 sky130_fd_sc_hd__nand2_1 _17498_ (.A(_01843_),
    .B(_01801_),
    .Y(_01844_));
 sky130_fd_sc_hd__mux2_1 _17499_ (.A0(\core.cpuregs[28][12] ),
    .A1(\core.cpuregs[29][12] ),
    .S(_01757_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _17500_ (.A0(\core.cpuregs[30][12] ),
    .A1(\core.cpuregs[31][12] ),
    .S(_01759_),
    .X(_01846_));
 sky130_fd_sc_hd__clkbuf_2 _17501_ (.A(_09617_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _17502_ (.A0(_01845_),
    .A1(_01846_),
    .S(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__nand2_1 _17503_ (.A(_01848_),
    .B(_01608_),
    .Y(_01849_));
 sky130_fd_sc_hd__mux2_1 _17504_ (.A0(\core.cpuregs[12][12] ),
    .A1(\core.cpuregs[13][12] ),
    .S(_01610_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _17505_ (.A0(\core.cpuregs[14][12] ),
    .A1(\core.cpuregs[15][12] ),
    .S(_10446_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _17506_ (.A0(_01850_),
    .A1(_01851_),
    .S(_01809_),
    .X(_01852_));
 sky130_fd_sc_hd__nand2_1 _17507_ (.A(_01852_),
    .B(_10449_),
    .Y(_01853_));
 sky130_fd_sc_hd__clkbuf_2 _17508_ (.A(_10371_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _17509_ (.A0(\core.cpuregs[8][12] ),
    .A1(\core.cpuregs[9][12] ),
    .S(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__clkbuf_2 _17510_ (.A(_04521_),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _17511_ (.A0(\core.cpuregs[10][12] ),
    .A1(\core.cpuregs[11][12] ),
    .S(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_2 _17512_ (.A0(_01855_),
    .A1(_01857_),
    .S(_01769_),
    .X(_01858_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_01858_),
    .B(_01618_),
    .Y(_01859_));
 sky130_fd_sc_hd__buf_1 _17514_ (.A(_10379_),
    .X(_01860_));
 sky130_fd_sc_hd__and3_1 _17515_ (.A(_01853_),
    .B(_01859_),
    .C(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__a31o_1 _17516_ (.A1(_01797_),
    .A2(_01844_),
    .A3(_01849_),
    .B1(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__a21oi_4 _17517_ (.A1(_01862_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01863_));
 sky130_fd_sc_hd__clkbuf_2 _17518_ (.A(_10339_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _17519_ (.A0(\core.cpuregs[16][12] ),
    .A1(\core.cpuregs[17][12] ),
    .S(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__clkbuf_2 _17520_ (.A(_10392_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _17521_ (.A0(\core.cpuregs[18][12] ),
    .A1(\core.cpuregs[19][12] ),
    .S(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _17522_ (.A0(_01865_),
    .A1(_01867_),
    .S(_01730_),
    .X(_01868_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17523_ (.A(_10399_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__clkbuf_2 _17525_ (.A(_10392_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _17526_ (.A0(\core.cpuregs[22][12] ),
    .A1(\core.cpuregs[23][12] ),
    .S(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__clkbuf_2 _17527_ (.A(_04522_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _17528_ (.A0(\core.cpuregs[20][12] ),
    .A1(\core.cpuregs[21][12] ),
    .S(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__clkbuf_2 _17529_ (.A(_04537_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _17530_ (.A0(_01872_),
    .A1(_01874_),
    .S(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_01876_),
    .B(_01630_),
    .Y(_01877_));
 sky130_fd_sc_hd__mux2_1 _17532_ (.A0(\core.cpuregs[6][12] ),
    .A1(\core.cpuregs[7][12] ),
    .S(_01783_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _17533_ (.A0(\core.cpuregs[4][12] ),
    .A1(\core.cpuregs[5][12] ),
    .S(_01785_),
    .X(_01879_));
 sky130_fd_sc_hd__clkbuf_2 _17534_ (.A(_09622_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _17535_ (.A0(_01878_),
    .A1(_01879_),
    .S(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__clkbuf_2 _17536_ (.A(_10418_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _17537_ (.A0(\core.cpuregs[0][12] ),
    .A1(\core.cpuregs[1][12] ),
    .S(_01637_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _17538_ (.A0(\core.cpuregs[2][12] ),
    .A1(\core.cpuregs[3][12] ),
    .S(_01639_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_2 _17539_ (.A0(_01883_),
    .A1(_01884_),
    .S(_01833_),
    .X(_01885_));
 sky130_fd_sc_hd__and2_1 _17540_ (.A(_01885_),
    .B(_01642_),
    .X(_01886_));
 sky130_fd_sc_hd__a211oi_1 _17541_ (.A1(_01633_),
    .A2(_01881_),
    .B1(_01882_),
    .C1(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a31o_1 _17542_ (.A1(_01819_),
    .A2(_01870_),
    .A3(_01877_),
    .B1(_01887_),
    .X(_01888_));
 sky130_fd_sc_hd__nand2_1 _17543_ (.A(_01888_),
    .B(_01747_),
    .Y(_01889_));
 sky130_fd_sc_hd__a22o_1 _17544_ (.A1(\core.decoded_imm[12] ),
    .A2(_10436_),
    .B1(_01863_),
    .B2(_01889_),
    .X(_01890_));
 sky130_fd_sc_hd__buf_4 _17545_ (.A(_10321_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _17546_ (.A0(_01890_),
    .A1(\core.pcpi_rs2[12] ),
    .S(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__clkbuf_1 _17547_ (.A(_01892_),
    .X(_00616_));
 sky130_fd_sc_hd__buf_2 _17548_ (.A(_04496_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _17549_ (.A0(\core.cpuregs[24][13] ),
    .A1(\core.cpuregs[25][13] ),
    .S(_01751_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _17550_ (.A0(\core.cpuregs[26][13] ),
    .A1(\core.cpuregs[27][13] ),
    .S(_01753_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_2 _17551_ (.A0(_01894_),
    .A1(_01895_),
    .S(_01708_),
    .X(_01896_));
 sky130_fd_sc_hd__nand2_8 _17552_ (.A(_01896_),
    .B(_01801_),
    .Y(_01897_));
 sky130_fd_sc_hd__mux2_1 _17553_ (.A0(\core.cpuregs[28][13] ),
    .A1(\core.cpuregs[29][13] ),
    .S(_01757_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _17554_ (.A0(\core.cpuregs[30][13] ),
    .A1(\core.cpuregs[31][13] ),
    .S(_01759_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_2 _17555_ (.A0(_01898_),
    .A1(_01899_),
    .S(_01847_),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_8 _17556_ (.A(_01900_),
    .B(_01608_),
    .Y(_01901_));
 sky130_fd_sc_hd__mux2_1 _17557_ (.A0(\core.cpuregs[12][13] ),
    .A1(\core.cpuregs[13][13] ),
    .S(_01610_),
    .X(_01902_));
 sky130_fd_sc_hd__clkbuf_2 _17558_ (.A(_10362_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _17559_ (.A0(\core.cpuregs[14][13] ),
    .A1(\core.cpuregs[15][13] ),
    .S(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _17560_ (.A0(_01902_),
    .A1(_01904_),
    .S(_01809_),
    .X(_01905_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17561_ (.A(_10368_),
    .X(_01906_));
 sky130_fd_sc_hd__nand2_1 _17562_ (.A(_01905_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__mux2_1 _17563_ (.A0(\core.cpuregs[8][13] ),
    .A1(\core.cpuregs[9][13] ),
    .S(_01854_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _17564_ (.A0(\core.cpuregs[10][13] ),
    .A1(\core.cpuregs[11][13] ),
    .S(_01856_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _17565_ (.A0(_01908_),
    .A1(_01909_),
    .S(_01769_),
    .X(_01910_));
 sky130_fd_sc_hd__nand2_1 _17566_ (.A(_01910_),
    .B(_01618_),
    .Y(_01911_));
 sky130_fd_sc_hd__and3_1 _17567_ (.A(_01907_),
    .B(_01911_),
    .C(_01860_),
    .X(_01912_));
 sky130_fd_sc_hd__a31o_1 _17568_ (.A1(_01797_),
    .A2(_01897_),
    .A3(_01901_),
    .B1(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__a21oi_2 _17569_ (.A1(_01913_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01914_));
 sky130_fd_sc_hd__mux2_1 _17570_ (.A0(\core.cpuregs[16][13] ),
    .A1(\core.cpuregs[17][13] ),
    .S(_01864_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _17571_ (.A0(\core.cpuregs[18][13] ),
    .A1(\core.cpuregs[19][13] ),
    .S(_01866_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _17572_ (.A0(_01915_),
    .A1(_01916_),
    .S(_01730_),
    .X(_01917_));
 sky130_fd_sc_hd__nand2_1 _17573_ (.A(_01917_),
    .B(_01869_),
    .Y(_01918_));
 sky130_fd_sc_hd__mux2_1 _17574_ (.A0(\core.cpuregs[22][13] ),
    .A1(\core.cpuregs[23][13] ),
    .S(_01871_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _17575_ (.A0(\core.cpuregs[20][13] ),
    .A1(\core.cpuregs[21][13] ),
    .S(_01873_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _17576_ (.A0(_01919_),
    .A1(_01920_),
    .S(_01875_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_1 _17577_ (.A(_01921_),
    .B(_01630_),
    .Y(_01922_));
 sky130_fd_sc_hd__mux2_1 _17578_ (.A0(\core.cpuregs[6][13] ),
    .A1(\core.cpuregs[7][13] ),
    .S(_01783_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _17579_ (.A0(\core.cpuregs[4][13] ),
    .A1(\core.cpuregs[5][13] ),
    .S(_01785_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _17580_ (.A0(_01923_),
    .A1(_01924_),
    .S(_01880_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _17581_ (.A0(\core.cpuregs[0][13] ),
    .A1(\core.cpuregs[1][13] ),
    .S(_01637_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _17582_ (.A0(\core.cpuregs[2][13] ),
    .A1(\core.cpuregs[3][13] ),
    .S(_01639_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _17583_ (.A0(_01926_),
    .A1(_01927_),
    .S(_01833_),
    .X(_01928_));
 sky130_fd_sc_hd__and2_1 _17584_ (.A(_01928_),
    .B(_01642_),
    .X(_01929_));
 sky130_fd_sc_hd__a211oi_1 _17585_ (.A1(_01633_),
    .A2(_01925_),
    .B1(_01882_),
    .C1(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__a31o_1 _17586_ (.A1(_01819_),
    .A2(_01918_),
    .A3(_01922_),
    .B1(_01930_),
    .X(_01931_));
 sky130_fd_sc_hd__nand2_1 _17587_ (.A(_01931_),
    .B(_01747_),
    .Y(_01932_));
 sky130_fd_sc_hd__a22o_1 _17588_ (.A1(\core.decoded_imm[13] ),
    .A2(_01893_),
    .B1(_01914_),
    .B2(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _17589_ (.A0(_01933_),
    .A1(\core.pcpi_rs2[13] ),
    .S(_01891_),
    .X(_01934_));
 sky130_fd_sc_hd__buf_1 _17590_ (.A(_01934_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _17591_ (.A0(\core.cpuregs[24][14] ),
    .A1(\core.cpuregs[25][14] ),
    .S(_01751_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _17592_ (.A0(\core.cpuregs[26][14] ),
    .A1(\core.cpuregs[27][14] ),
    .S(_01753_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _17593_ (.A0(_01935_),
    .A1(_01936_),
    .S(_01708_),
    .X(_01937_));
 sky130_fd_sc_hd__nand2_1 _17594_ (.A(_01937_),
    .B(_01801_),
    .Y(_01938_));
 sky130_fd_sc_hd__mux2_4 _17595_ (.A0(\core.cpuregs[28][14] ),
    .A1(\core.cpuregs[29][14] ),
    .S(_01757_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _17596_ (.A0(\core.cpuregs[30][14] ),
    .A1(\core.cpuregs[31][14] ),
    .S(_01759_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _17597_ (.A0(_01939_),
    .A1(_01940_),
    .S(_01847_),
    .X(_01941_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17598_ (.A(_10357_),
    .X(_01942_));
 sky130_fd_sc_hd__nand2_1 _17599_ (.A(_01941_),
    .B(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__clkbuf_2 _17600_ (.A(_10362_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _17601_ (.A0(\core.cpuregs[12][14] ),
    .A1(\core.cpuregs[13][14] ),
    .S(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _17602_ (.A0(\core.cpuregs[14][14] ),
    .A1(\core.cpuregs[15][14] ),
    .S(_01903_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _17603_ (.A0(_01945_),
    .A1(_01946_),
    .S(_01809_),
    .X(_01947_));
 sky130_fd_sc_hd__nand2_1 _17604_ (.A(_01947_),
    .B(_01906_),
    .Y(_01948_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(\core.cpuregs[8][14] ),
    .A1(\core.cpuregs[9][14] ),
    .S(_01854_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _17606_ (.A0(\core.cpuregs[10][14] ),
    .A1(\core.cpuregs[11][14] ),
    .S(_01856_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _17607_ (.A0(_01949_),
    .A1(_01950_),
    .S(_01769_),
    .X(_01951_));
 sky130_fd_sc_hd__clkbuf_4 _17608_ (.A(_10346_),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _17609_ (.A(_01951_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__and3_1 _17610_ (.A(_01948_),
    .B(_01953_),
    .C(_01860_),
    .X(_01954_));
 sky130_fd_sc_hd__a31o_1 _17611_ (.A1(_01797_),
    .A2(_01938_),
    .A3(_01943_),
    .B1(_01954_),
    .X(_01955_));
 sky130_fd_sc_hd__a21oi_1 _17612_ (.A1(_01955_),
    .A2(_01725_),
    .B1(_01726_),
    .Y(_01956_));
 sky130_fd_sc_hd__mux2_1 _17613_ (.A0(\core.cpuregs[16][14] ),
    .A1(\core.cpuregs[17][14] ),
    .S(_01864_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _17614_ (.A0(\core.cpuregs[18][14] ),
    .A1(\core.cpuregs[19][14] ),
    .S(_01866_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_8 _17615_ (.A0(_01957_),
    .A1(_01958_),
    .S(_01730_),
    .X(_01959_));
 sky130_fd_sc_hd__nand2_1 _17616_ (.A(_01959_),
    .B(_01869_),
    .Y(_01960_));
 sky130_fd_sc_hd__mux2_2 _17617_ (.A0(\core.cpuregs[22][14] ),
    .A1(\core.cpuregs[23][14] ),
    .S(_01871_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _17618_ (.A0(\core.cpuregs[20][14] ),
    .A1(\core.cpuregs[21][14] ),
    .S(_01873_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _17619_ (.A0(_01961_),
    .A1(_01962_),
    .S(_01875_),
    .X(_01963_));
 sky130_fd_sc_hd__buf_2 _17620_ (.A(_10369_),
    .X(_01964_));
 sky130_fd_sc_hd__nand2_1 _17621_ (.A(_01963_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__clkbuf_2 _17622_ (.A(_10357_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _17623_ (.A0(\core.cpuregs[6][14] ),
    .A1(\core.cpuregs[7][14] ),
    .S(_01783_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _17624_ (.A0(\core.cpuregs[4][14] ),
    .A1(\core.cpuregs[5][14] ),
    .S(_01785_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _17625_ (.A0(_01967_),
    .A1(_01968_),
    .S(_01880_),
    .X(_01969_));
 sky130_fd_sc_hd__buf_4 _17626_ (.A(_09648_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _17627_ (.A0(\core.cpuregs[0][14] ),
    .A1(\core.cpuregs[1][14] ),
    .S(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__clkbuf_2 _17628_ (.A(_10338_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _17629_ (.A0(\core.cpuregs[2][14] ),
    .A1(\core.cpuregs[3][14] ),
    .S(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _17630_ (.A0(_01971_),
    .A1(_01973_),
    .S(_01833_),
    .X(_01974_));
 sky130_fd_sc_hd__clkbuf_4 _17631_ (.A(_10346_),
    .X(_01975_));
 sky130_fd_sc_hd__and2_1 _17632_ (.A(_01974_),
    .B(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__a211oi_2 _17633_ (.A1(_01966_),
    .A2(_01969_),
    .B1(_01882_),
    .C1(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__a31o_4 _17634_ (.A1(_01819_),
    .A2(_01960_),
    .A3(_01965_),
    .B1(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__nand2_1 _17635_ (.A(_01978_),
    .B(_01747_),
    .Y(_01979_));
 sky130_fd_sc_hd__a22o_1 _17636_ (.A1(\core.decoded_imm[14] ),
    .A2(_01893_),
    .B1(_01956_),
    .B2(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _17637_ (.A0(_01980_),
    .A1(\core.pcpi_rs2[14] ),
    .S(_01891_),
    .X(_01981_));
 sky130_fd_sc_hd__clkbuf_1 _17638_ (.A(_01981_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _17639_ (.A0(\core.cpuregs[24][15] ),
    .A1(\core.cpuregs[25][15] ),
    .S(_01751_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _17640_ (.A0(\core.cpuregs[26][15] ),
    .A1(\core.cpuregs[27][15] ),
    .S(_01753_),
    .X(_01983_));
 sky130_fd_sc_hd__clkbuf_2 _17641_ (.A(_04641_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_2 _17642_ (.A0(_01982_),
    .A1(_01983_),
    .S(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__nand2_8 _17643_ (.A(_01985_),
    .B(_01801_),
    .Y(_01986_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(\core.cpuregs[28][15] ),
    .A1(\core.cpuregs[29][15] ),
    .S(_01757_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_2 _17645_ (.A0(\core.cpuregs[30][15] ),
    .A1(\core.cpuregs[31][15] ),
    .S(_01759_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _17646_ (.A0(_01987_),
    .A1(_01988_),
    .S(_01847_),
    .X(_01989_));
 sky130_fd_sc_hd__nand2_1 _17647_ (.A(_01989_),
    .B(_01942_),
    .Y(_01990_));
 sky130_fd_sc_hd__mux2_1 _17648_ (.A0(\core.cpuregs[12][15] ),
    .A1(\core.cpuregs[13][15] ),
    .S(_01944_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _17649_ (.A0(\core.cpuregs[14][15] ),
    .A1(\core.cpuregs[15][15] ),
    .S(_01903_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(_01991_),
    .A1(_01992_),
    .S(_01809_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _17651_ (.A(_01993_),
    .B(_01906_),
    .Y(_01994_));
 sky130_fd_sc_hd__mux2_1 _17652_ (.A0(\core.cpuregs[8][15] ),
    .A1(\core.cpuregs[9][15] ),
    .S(_01854_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _17653_ (.A0(\core.cpuregs[10][15] ),
    .A1(\core.cpuregs[11][15] ),
    .S(_01856_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_8 _17654_ (.A0(_01995_),
    .A1(_01996_),
    .S(_01769_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_01997_),
    .B(_01952_),
    .Y(_01998_));
 sky130_fd_sc_hd__and3_1 _17656_ (.A(_01994_),
    .B(_01998_),
    .C(_01860_),
    .X(_01999_));
 sky130_fd_sc_hd__a31o_2 _17657_ (.A1(_01797_),
    .A2(_01986_),
    .A3(_01990_),
    .B1(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__clkbuf_4 _17658_ (.A(_10383_),
    .X(_02001_));
 sky130_fd_sc_hd__clkbuf_4 _17659_ (.A(_10386_),
    .X(_02002_));
 sky130_fd_sc_hd__a21oi_1 _17660_ (.A1(_02000_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__mux2_8 _17661_ (.A0(\core.cpuregs[16][15] ),
    .A1(\core.cpuregs[17][15] ),
    .S(_01864_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _17662_ (.A0(\core.cpuregs[18][15] ),
    .A1(\core.cpuregs[19][15] ),
    .S(_01866_),
    .X(_02005_));
 sky130_fd_sc_hd__clkbuf_2 _17663_ (.A(_10395_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _17664_ (.A0(_02004_),
    .A1(_02005_),
    .S(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__nand2_1 _17665_ (.A(_02007_),
    .B(_01869_),
    .Y(_02008_));
 sky130_fd_sc_hd__mux2_1 _17666_ (.A0(\core.cpuregs[22][15] ),
    .A1(\core.cpuregs[23][15] ),
    .S(_01871_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _17667_ (.A0(\core.cpuregs[20][15] ),
    .A1(\core.cpuregs[21][15] ),
    .S(_01873_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _17668_ (.A0(_02009_),
    .A1(_02010_),
    .S(_01875_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(_02011_),
    .B(_01964_),
    .Y(_02012_));
 sky130_fd_sc_hd__mux2_1 _17670_ (.A0(\core.cpuregs[6][15] ),
    .A1(\core.cpuregs[7][15] ),
    .S(_01783_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _17671_ (.A0(\core.cpuregs[4][15] ),
    .A1(\core.cpuregs[5][15] ),
    .S(_01785_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _17672_ (.A0(_02013_),
    .A1(_02014_),
    .S(_01880_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(\core.cpuregs[0][15] ),
    .A1(\core.cpuregs[1][15] ),
    .S(_01970_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _17674_ (.A0(\core.cpuregs[2][15] ),
    .A1(\core.cpuregs[3][15] ),
    .S(_01972_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(_02016_),
    .A1(_02017_),
    .S(_01833_),
    .X(_02018_));
 sky130_fd_sc_hd__and2_1 _17676_ (.A(_02018_),
    .B(_01975_),
    .X(_02019_));
 sky130_fd_sc_hd__a211oi_2 _17677_ (.A1(_01966_),
    .A2(_02015_),
    .B1(_01882_),
    .C1(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__a31o_4 _17678_ (.A1(_01819_),
    .A2(_02008_),
    .A3(_02012_),
    .B1(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_2 _17679_ (.A(_01746_),
    .X(_02022_));
 sky130_fd_sc_hd__nand2_1 _17680_ (.A(_02021_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__a22o_1 _17681_ (.A1(\core.decoded_imm[15] ),
    .A2(_01893_),
    .B1(_02003_),
    .B2(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _17682_ (.A0(_02024_),
    .A1(\core.pcpi_rs2[15] ),
    .S(_01891_),
    .X(_02025_));
 sky130_fd_sc_hd__buf_1 _17683_ (.A(_02025_),
    .X(_00619_));
 sky130_fd_sc_hd__clkbuf_2 _17684_ (.A(_04567_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(\core.cpuregs[24][16] ),
    .A1(\core.cpuregs[25][16] ),
    .S(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__clkbuf_2 _17686_ (.A(_04636_),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _17687_ (.A0(\core.cpuregs[26][16] ),
    .A1(\core.cpuregs[27][16] ),
    .S(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__mux2_1 _17688_ (.A0(_02027_),
    .A1(_02029_),
    .S(_01984_),
    .X(_02030_));
 sky130_fd_sc_hd__nand2_1 _17689_ (.A(_02030_),
    .B(_01801_),
    .Y(_02031_));
 sky130_fd_sc_hd__clkbuf_2 _17690_ (.A(_04662_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _17691_ (.A0(\core.cpuregs[28][16] ),
    .A1(\core.cpuregs[29][16] ),
    .S(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__clkbuf_2 _17692_ (.A(_10352_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(\core.cpuregs[30][16] ),
    .A1(\core.cpuregs[31][16] ),
    .S(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_8 _17694_ (.A0(_02033_),
    .A1(_02035_),
    .S(_01847_),
    .X(_02036_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(_02036_),
    .B(_01942_),
    .Y(_02037_));
 sky130_fd_sc_hd__mux2_1 _17696_ (.A0(\core.cpuregs[12][16] ),
    .A1(\core.cpuregs[13][16] ),
    .S(_01944_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _17697_ (.A0(\core.cpuregs[14][16] ),
    .A1(\core.cpuregs[15][16] ),
    .S(_01903_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(_02038_),
    .A1(_02039_),
    .S(_01809_),
    .X(_02040_));
 sky130_fd_sc_hd__nand2_1 _17699_ (.A(_02040_),
    .B(_01906_),
    .Y(_02041_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(\core.cpuregs[8][16] ),
    .A1(\core.cpuregs[9][16] ),
    .S(_01854_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _17701_ (.A0(\core.cpuregs[10][16] ),
    .A1(\core.cpuregs[11][16] ),
    .S(_01856_),
    .X(_02043_));
 sky130_fd_sc_hd__clkbuf_2 _17702_ (.A(_04640_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _17703_ (.A0(_02042_),
    .A1(_02043_),
    .S(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_1 _17704_ (.A(_02045_),
    .B(_01952_),
    .Y(_02046_));
 sky130_fd_sc_hd__and3_2 _17705_ (.A(_02041_),
    .B(_02046_),
    .C(_01860_),
    .X(_02047_));
 sky130_fd_sc_hd__a31o_2 _17706_ (.A1(_01797_),
    .A2(_02031_),
    .A3(_02037_),
    .B1(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__a21oi_4 _17707_ (.A1(_02048_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02049_));
 sky130_fd_sc_hd__mux2_1 _17708_ (.A0(\core.cpuregs[16][16] ),
    .A1(\core.cpuregs[17][16] ),
    .S(_01864_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _17709_ (.A0(\core.cpuregs[18][16] ),
    .A1(\core.cpuregs[19][16] ),
    .S(_01866_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _17710_ (.A0(_02050_),
    .A1(_02051_),
    .S(_02006_),
    .X(_02052_));
 sky130_fd_sc_hd__nand2_1 _17711_ (.A(_02052_),
    .B(_01869_),
    .Y(_02053_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(\core.cpuregs[22][16] ),
    .A1(\core.cpuregs[23][16] ),
    .S(_01871_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _17713_ (.A0(\core.cpuregs[20][16] ),
    .A1(\core.cpuregs[21][16] ),
    .S(_01873_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_2 _17714_ (.A0(_02054_),
    .A1(_02055_),
    .S(_01875_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_8 _17715_ (.A(_02056_),
    .B(_01964_),
    .Y(_02057_));
 sky130_fd_sc_hd__clkbuf_4 _17716_ (.A(_10413_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _17717_ (.A0(\core.cpuregs[6][16] ),
    .A1(\core.cpuregs[7][16] ),
    .S(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__clkbuf_4 _17718_ (.A(_10413_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _17719_ (.A0(\core.cpuregs[4][16] ),
    .A1(\core.cpuregs[5][16] ),
    .S(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _17720_ (.A0(_02059_),
    .A1(_02061_),
    .S(_01880_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _17721_ (.A0(\core.cpuregs[0][16] ),
    .A1(\core.cpuregs[1][16] ),
    .S(_01970_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _17722_ (.A0(\core.cpuregs[2][16] ),
    .A1(\core.cpuregs[3][16] ),
    .S(_01972_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _17723_ (.A0(_02063_),
    .A1(_02064_),
    .S(_01833_),
    .X(_02065_));
 sky130_fd_sc_hd__and2_2 _17724_ (.A(_02065_),
    .B(_01975_),
    .X(_02066_));
 sky130_fd_sc_hd__a211oi_2 _17725_ (.A1(_01966_),
    .A2(_02062_),
    .B1(_01882_),
    .C1(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__a31o_1 _17726_ (.A1(_01819_),
    .A2(_02053_),
    .A3(_02057_),
    .B1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nand2_1 _17727_ (.A(_02068_),
    .B(_02022_),
    .Y(_02069_));
 sky130_fd_sc_hd__a22o_1 _17728_ (.A1(\core.decoded_imm[16] ),
    .A2(_01893_),
    .B1(_02049_),
    .B2(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _17729_ (.A0(_02070_),
    .A1(\core.pcpi_rs2[16] ),
    .S(_01891_),
    .X(_02071_));
 sky130_fd_sc_hd__clkbuf_1 _17730_ (.A(_02071_),
    .X(_00620_));
 sky130_fd_sc_hd__buf_2 _17731_ (.A(_10418_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _17732_ (.A0(\core.cpuregs[24][17] ),
    .A1(\core.cpuregs[25][17] ),
    .S(_02026_),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_1 _17733_ (.A0(\core.cpuregs[26][17] ),
    .A1(\core.cpuregs[27][17] ),
    .S(_02028_),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _17734_ (.A0(_02073_),
    .A1(_02074_),
    .S(_01984_),
    .X(_02075_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17735_ (.A(_10347_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_02075_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__mux2_1 _17737_ (.A0(\core.cpuregs[28][17] ),
    .A1(\core.cpuregs[29][17] ),
    .S(_02032_),
    .X(_02078_));
 sky130_fd_sc_hd__mux2_1 _17738_ (.A0(\core.cpuregs[30][17] ),
    .A1(\core.cpuregs[31][17] ),
    .S(_02034_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_1 _17739_ (.A0(_02078_),
    .A1(_02079_),
    .S(_01847_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_1 _17740_ (.A(_02080_),
    .B(_01942_),
    .Y(_02081_));
 sky130_fd_sc_hd__mux2_1 _17741_ (.A0(\core.cpuregs[12][17] ),
    .A1(\core.cpuregs[13][17] ),
    .S(_01944_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _17742_ (.A0(\core.cpuregs[14][17] ),
    .A1(\core.cpuregs[15][17] ),
    .S(_01903_),
    .X(_02083_));
 sky130_fd_sc_hd__clkbuf_4 _17743_ (.A(_10365_),
    .X(_02084_));
 sky130_fd_sc_hd__mux2_1 _17744_ (.A0(_02082_),
    .A1(_02083_),
    .S(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _17745_ (.A(_02085_),
    .B(_01906_),
    .Y(_02086_));
 sky130_fd_sc_hd__mux2_1 _17746_ (.A0(\core.cpuregs[8][17] ),
    .A1(\core.cpuregs[9][17] ),
    .S(_01854_),
    .X(_02087_));
 sky130_fd_sc_hd__mux2_1 _17747_ (.A0(\core.cpuregs[10][17] ),
    .A1(\core.cpuregs[11][17] ),
    .S(_01856_),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _17748_ (.A0(_02087_),
    .A1(_02088_),
    .S(_02044_),
    .X(_02089_));
 sky130_fd_sc_hd__nand2_1 _17749_ (.A(_02089_),
    .B(_01952_),
    .Y(_02090_));
 sky130_fd_sc_hd__and3_1 _17750_ (.A(_02086_),
    .B(_02090_),
    .C(_01860_),
    .X(_02091_));
 sky130_fd_sc_hd__a31o_2 _17751_ (.A1(_02072_),
    .A2(_02077_),
    .A3(_02081_),
    .B1(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__a21oi_4 _17752_ (.A1(_02092_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02093_));
 sky130_fd_sc_hd__clkbuf_4 _17753_ (.A(_10336_),
    .X(_02094_));
 sky130_fd_sc_hd__mux2_1 _17754_ (.A0(\core.cpuregs[16][17] ),
    .A1(\core.cpuregs[17][17] ),
    .S(_01864_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _17755_ (.A0(\core.cpuregs[18][17] ),
    .A1(\core.cpuregs[19][17] ),
    .S(_01866_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _17756_ (.A0(_02095_),
    .A1(_02096_),
    .S(_02006_),
    .X(_02097_));
 sky130_fd_sc_hd__nand2_1 _17757_ (.A(_02097_),
    .B(_01869_),
    .Y(_02098_));
 sky130_fd_sc_hd__mux2_1 _17758_ (.A0(\core.cpuregs[22][17] ),
    .A1(\core.cpuregs[23][17] ),
    .S(_01871_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _17759_ (.A0(\core.cpuregs[20][17] ),
    .A1(\core.cpuregs[21][17] ),
    .S(_01873_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_2 _17760_ (.A0(_02099_),
    .A1(_02100_),
    .S(_01875_),
    .X(_02101_));
 sky130_fd_sc_hd__nand2_1 _17761_ (.A(_02101_),
    .B(_01964_),
    .Y(_02102_));
 sky130_fd_sc_hd__mux2_1 _17762_ (.A0(\core.cpuregs[6][17] ),
    .A1(\core.cpuregs[7][17] ),
    .S(_02058_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _17763_ (.A0(\core.cpuregs[4][17] ),
    .A1(\core.cpuregs[5][17] ),
    .S(_02060_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _17764_ (.A0(_02103_),
    .A1(_02104_),
    .S(_01880_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _17765_ (.A0(\core.cpuregs[0][17] ),
    .A1(\core.cpuregs[1][17] ),
    .S(_01970_),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _17766_ (.A0(\core.cpuregs[2][17] ),
    .A1(\core.cpuregs[3][17] ),
    .S(_01972_),
    .X(_02107_));
 sky130_fd_sc_hd__clkbuf_4 _17767_ (.A(_09650_),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _17768_ (.A0(_02106_),
    .A1(_02107_),
    .S(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__and2_1 _17769_ (.A(_02109_),
    .B(_01975_),
    .X(_02110_));
 sky130_fd_sc_hd__a211oi_2 _17770_ (.A1(_01966_),
    .A2(_02105_),
    .B1(_01882_),
    .C1(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__a31o_1 _17771_ (.A1(_02094_),
    .A2(_02098_),
    .A3(_02102_),
    .B1(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _17772_ (.A(_02112_),
    .B(_02022_),
    .Y(_02113_));
 sky130_fd_sc_hd__a22o_1 _17773_ (.A1(\core.decoded_imm[17] ),
    .A2(_01893_),
    .B1(_02093_),
    .B2(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _17774_ (.A0(_02114_),
    .A1(\core.pcpi_rs2[17] ),
    .S(_01891_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_1 _17775_ (.A(_02115_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _17776_ (.A0(\core.cpuregs[24][18] ),
    .A1(\core.cpuregs[25][18] ),
    .S(_02026_),
    .X(_02116_));
 sky130_fd_sc_hd__mux2_1 _17777_ (.A0(\core.cpuregs[26][18] ),
    .A1(\core.cpuregs[27][18] ),
    .S(_02028_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _17778_ (.A0(_02116_),
    .A1(_02117_),
    .S(_01984_),
    .X(_02118_));
 sky130_fd_sc_hd__nand2_1 _17779_ (.A(_02118_),
    .B(_02076_),
    .Y(_02119_));
 sky130_fd_sc_hd__mux2_1 _17780_ (.A0(\core.cpuregs[28][18] ),
    .A1(\core.cpuregs[29][18] ),
    .S(_02032_),
    .X(_02120_));
 sky130_fd_sc_hd__mux2_1 _17781_ (.A0(\core.cpuregs[30][18] ),
    .A1(\core.cpuregs[31][18] ),
    .S(_02034_),
    .X(_02121_));
 sky130_fd_sc_hd__clkbuf_2 _17782_ (.A(_09617_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _17783_ (.A0(_02120_),
    .A1(_02121_),
    .S(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__nand2_1 _17784_ (.A(_02123_),
    .B(_01942_),
    .Y(_02124_));
 sky130_fd_sc_hd__mux2_1 _17785_ (.A0(\core.cpuregs[12][18] ),
    .A1(\core.cpuregs[13][18] ),
    .S(_01944_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _17786_ (.A0(\core.cpuregs[14][18] ),
    .A1(\core.cpuregs[15][18] ),
    .S(_01903_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _17787_ (.A0(_02125_),
    .A1(_02126_),
    .S(_02084_),
    .X(_02127_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_02127_),
    .B(_01906_),
    .Y(_02128_));
 sky130_fd_sc_hd__clkbuf_4 _17789_ (.A(_10371_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _17790_ (.A0(\core.cpuregs[8][18] ),
    .A1(\core.cpuregs[9][18] ),
    .S(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__clkbuf_4 _17791_ (.A(_04521_),
    .X(_02131_));
 sky130_fd_sc_hd__mux2_1 _17792_ (.A0(\core.cpuregs[10][18] ),
    .A1(\core.cpuregs[11][18] ),
    .S(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_2 _17793_ (.A0(_02130_),
    .A1(_02132_),
    .S(_02044_),
    .X(_02133_));
 sky130_fd_sc_hd__nand2_1 _17794_ (.A(_02133_),
    .B(_01952_),
    .Y(_02134_));
 sky130_fd_sc_hd__clkbuf_4 _17795_ (.A(_10379_),
    .X(_02135_));
 sky130_fd_sc_hd__and3_1 _17796_ (.A(_02128_),
    .B(_02134_),
    .C(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__a31o_1 _17797_ (.A1(_02072_),
    .A2(_02119_),
    .A3(_02124_),
    .B1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__a21oi_1 _17798_ (.A1(_02137_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02138_));
 sky130_fd_sc_hd__buf_4 _17799_ (.A(_10339_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_4 _17800_ (.A0(\core.cpuregs[16][18] ),
    .A1(\core.cpuregs[17][18] ),
    .S(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_2 _17801_ (.A(_10392_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _17802_ (.A0(\core.cpuregs[18][18] ),
    .A1(\core.cpuregs[19][18] ),
    .S(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _17803_ (.A0(_02140_),
    .A1(_02142_),
    .S(_02006_),
    .X(_02143_));
 sky130_fd_sc_hd__clkbuf_2 _17804_ (.A(_10399_),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _17805_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__buf_4 _17806_ (.A(_04522_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _17807_ (.A0(\core.cpuregs[22][18] ),
    .A1(\core.cpuregs[23][18] ),
    .S(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__buf_4 _17808_ (.A(_04532_),
    .X(_02148_));
 sky130_fd_sc_hd__mux2_1 _17809_ (.A0(\core.cpuregs[20][18] ),
    .A1(\core.cpuregs[21][18] ),
    .S(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__clkbuf_4 _17810_ (.A(_04537_),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _17811_ (.A0(_02147_),
    .A1(_02149_),
    .S(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__nand2_1 _17812_ (.A(_02151_),
    .B(_01964_),
    .Y(_02152_));
 sky130_fd_sc_hd__mux2_1 _17813_ (.A0(\core.cpuregs[6][18] ),
    .A1(\core.cpuregs[7][18] ),
    .S(_02058_),
    .X(_02153_));
 sky130_fd_sc_hd__mux2_1 _17814_ (.A0(\core.cpuregs[4][18] ),
    .A1(\core.cpuregs[5][18] ),
    .S(_02060_),
    .X(_02154_));
 sky130_fd_sc_hd__clkbuf_2 _17815_ (.A(_09622_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _17816_ (.A0(_02153_),
    .A1(_02154_),
    .S(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__clkbuf_2 _17817_ (.A(_10418_),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _17818_ (.A0(\core.cpuregs[0][18] ),
    .A1(\core.cpuregs[1][18] ),
    .S(_01970_),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _17819_ (.A0(\core.cpuregs[2][18] ),
    .A1(\core.cpuregs[3][18] ),
    .S(_01972_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _17820_ (.A0(_02158_),
    .A1(_02159_),
    .S(_02108_),
    .X(_02160_));
 sky130_fd_sc_hd__and2_1 _17821_ (.A(_02160_),
    .B(_01975_),
    .X(_02161_));
 sky130_fd_sc_hd__a211oi_2 _17822_ (.A1(_01966_),
    .A2(_02156_),
    .B1(_02157_),
    .C1(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__a31o_1 _17823_ (.A1(_02094_),
    .A2(_02145_),
    .A3(_02152_),
    .B1(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__nand2_2 _17824_ (.A(_02163_),
    .B(_02022_),
    .Y(_02164_));
 sky130_fd_sc_hd__a22o_1 _17825_ (.A1(\core.decoded_imm[18] ),
    .A2(_01893_),
    .B1(_02138_),
    .B2(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__buf_2 _17826_ (.A(_10321_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _17827_ (.A0(_02165_),
    .A1(\core.pcpi_rs2[18] ),
    .S(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17828_ (.A(_02167_),
    .X(_00622_));
 sky130_fd_sc_hd__buf_2 _17829_ (.A(_04496_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _17830_ (.A0(\core.cpuregs[24][19] ),
    .A1(\core.cpuregs[25][19] ),
    .S(_02026_),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_1 _17831_ (.A0(\core.cpuregs[26][19] ),
    .A1(\core.cpuregs[27][19] ),
    .S(_02028_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _17832_ (.A0(_02169_),
    .A1(_02170_),
    .S(_01984_),
    .X(_02171_));
 sky130_fd_sc_hd__nand2_1 _17833_ (.A(_02171_),
    .B(_02076_),
    .Y(_02172_));
 sky130_fd_sc_hd__mux2_1 _17834_ (.A0(\core.cpuregs[28][19] ),
    .A1(\core.cpuregs[29][19] ),
    .S(_02032_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _17835_ (.A0(\core.cpuregs[30][19] ),
    .A1(\core.cpuregs[31][19] ),
    .S(_02034_),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_2 _17836_ (.A0(_02173_),
    .A1(_02174_),
    .S(_02122_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2_1 _17837_ (.A(_02175_),
    .B(_01942_),
    .Y(_02176_));
 sky130_fd_sc_hd__mux2_1 _17838_ (.A0(\core.cpuregs[12][19] ),
    .A1(\core.cpuregs[13][19] ),
    .S(_01944_),
    .X(_02177_));
 sky130_fd_sc_hd__clkbuf_4 _17839_ (.A(_10371_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _17840_ (.A0(\core.cpuregs[14][19] ),
    .A1(\core.cpuregs[15][19] ),
    .S(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _17841_ (.A0(_02177_),
    .A1(_02179_),
    .S(_02084_),
    .X(_02180_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17842_ (.A(_10368_),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_1 _17843_ (.A(_02180_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__mux2_1 _17844_ (.A0(\core.cpuregs[8][19] ),
    .A1(\core.cpuregs[9][19] ),
    .S(_02129_),
    .X(_02183_));
 sky130_fd_sc_hd__mux2_1 _17845_ (.A0(\core.cpuregs[10][19] ),
    .A1(\core.cpuregs[11][19] ),
    .S(_02131_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _17846_ (.A0(_02183_),
    .A1(_02184_),
    .S(_02044_),
    .X(_02185_));
 sky130_fd_sc_hd__nand2_1 _17847_ (.A(_02185_),
    .B(_01952_),
    .Y(_02186_));
 sky130_fd_sc_hd__and3_1 _17848_ (.A(_02182_),
    .B(_02186_),
    .C(_02135_),
    .X(_02187_));
 sky130_fd_sc_hd__a31o_1 _17849_ (.A1(_02072_),
    .A2(_02172_),
    .A3(_02176_),
    .B1(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__a21oi_1 _17850_ (.A1(_02188_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02189_));
 sky130_fd_sc_hd__mux2_1 _17851_ (.A0(\core.cpuregs[16][19] ),
    .A1(\core.cpuregs[17][19] ),
    .S(_02139_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _17852_ (.A0(\core.cpuregs[18][19] ),
    .A1(\core.cpuregs[19][19] ),
    .S(_02141_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _17853_ (.A0(_02190_),
    .A1(_02191_),
    .S(_02006_),
    .X(_02192_));
 sky130_fd_sc_hd__nand2_1 _17854_ (.A(_02192_),
    .B(_02144_),
    .Y(_02193_));
 sky130_fd_sc_hd__mux2_1 _17855_ (.A0(\core.cpuregs[22][19] ),
    .A1(\core.cpuregs[23][19] ),
    .S(_02146_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _17856_ (.A0(\core.cpuregs[20][19] ),
    .A1(\core.cpuregs[21][19] ),
    .S(_02148_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _17857_ (.A0(_02194_),
    .A1(_02195_),
    .S(_02150_),
    .X(_02196_));
 sky130_fd_sc_hd__nand2_1 _17858_ (.A(_02196_),
    .B(_01964_),
    .Y(_02197_));
 sky130_fd_sc_hd__mux2_1 _17859_ (.A0(\core.cpuregs[6][19] ),
    .A1(\core.cpuregs[7][19] ),
    .S(_02058_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _17860_ (.A0(\core.cpuregs[4][19] ),
    .A1(\core.cpuregs[5][19] ),
    .S(_02060_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_2 _17861_ (.A0(_02198_),
    .A1(_02199_),
    .S(_02155_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _17862_ (.A0(\core.cpuregs[0][19] ),
    .A1(\core.cpuregs[1][19] ),
    .S(_01970_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _17863_ (.A0(\core.cpuregs[2][19] ),
    .A1(\core.cpuregs[3][19] ),
    .S(_01972_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _17864_ (.A0(_02201_),
    .A1(_02202_),
    .S(_02108_),
    .X(_02203_));
 sky130_fd_sc_hd__and2_1 _17865_ (.A(_02203_),
    .B(_01975_),
    .X(_02204_));
 sky130_fd_sc_hd__a211oi_1 _17866_ (.A1(_01966_),
    .A2(_02200_),
    .B1(_02157_),
    .C1(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__a31o_1 _17867_ (.A1(_02094_),
    .A2(_02193_),
    .A3(_02197_),
    .B1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__nand2_2 _17868_ (.A(_02206_),
    .B(_02022_),
    .Y(_02207_));
 sky130_fd_sc_hd__a22o_1 _17869_ (.A1(\core.decoded_imm[19] ),
    .A2(_02168_),
    .B1(_02189_),
    .B2(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_2 _17870_ (.A0(_02208_),
    .A1(\core.pcpi_rs2[19] ),
    .S(_02166_),
    .X(_02209_));
 sky130_fd_sc_hd__clkbuf_1 _17871_ (.A(_02209_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _17872_ (.A0(\core.cpuregs[24][20] ),
    .A1(\core.cpuregs[25][20] ),
    .S(_02026_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _17873_ (.A0(\core.cpuregs[26][20] ),
    .A1(\core.cpuregs[27][20] ),
    .S(_02028_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _17874_ (.A0(_02210_),
    .A1(_02211_),
    .S(_01984_),
    .X(_02212_));
 sky130_fd_sc_hd__nand2_1 _17875_ (.A(_02212_),
    .B(_02076_),
    .Y(_02213_));
 sky130_fd_sc_hd__mux2_1 _17876_ (.A0(\core.cpuregs[28][20] ),
    .A1(\core.cpuregs[29][20] ),
    .S(_02032_),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _17877_ (.A0(\core.cpuregs[30][20] ),
    .A1(\core.cpuregs[31][20] ),
    .S(_02034_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _17878_ (.A0(_02214_),
    .A1(_02215_),
    .S(_02122_),
    .X(_02216_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17879_ (.A(_10368_),
    .X(_02217_));
 sky130_fd_sc_hd__nand2_1 _17880_ (.A(_02216_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__clkbuf_4 _17881_ (.A(_10362_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _17882_ (.A0(\core.cpuregs[12][20] ),
    .A1(\core.cpuregs[13][20] ),
    .S(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _17883_ (.A0(\core.cpuregs[14][20] ),
    .A1(\core.cpuregs[15][20] ),
    .S(_02178_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _17884_ (.A0(_02220_),
    .A1(_02221_),
    .S(_02084_),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_1 _17885_ (.A(_02222_),
    .B(_02181_),
    .Y(_02223_));
 sky130_fd_sc_hd__mux2_1 _17886_ (.A0(\core.cpuregs[8][20] ),
    .A1(\core.cpuregs[9][20] ),
    .S(_02129_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _17887_ (.A0(\core.cpuregs[10][20] ),
    .A1(\core.cpuregs[11][20] ),
    .S(_02131_),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _17888_ (.A0(_02224_),
    .A1(_02225_),
    .S(_02044_),
    .X(_02226_));
 sky130_fd_sc_hd__clkbuf_4 _17889_ (.A(_10346_),
    .X(_02227_));
 sky130_fd_sc_hd__nand2_1 _17890_ (.A(_02226_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__and3_1 _17891_ (.A(_02223_),
    .B(_02228_),
    .C(_02135_),
    .X(_02229_));
 sky130_fd_sc_hd__a31o_1 _17892_ (.A1(_02072_),
    .A2(_02213_),
    .A3(_02218_),
    .B1(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__a21oi_4 _17893_ (.A1(_02230_),
    .A2(_02001_),
    .B1(_02002_),
    .Y(_02231_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(\core.cpuregs[16][20] ),
    .A1(\core.cpuregs[17][20] ),
    .S(_02139_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_2 _17895_ (.A0(\core.cpuregs[18][20] ),
    .A1(\core.cpuregs[19][20] ),
    .S(_02141_),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _17896_ (.A0(_02232_),
    .A1(_02233_),
    .S(_02006_),
    .X(_02234_));
 sky130_fd_sc_hd__nand2_1 _17897_ (.A(_02234_),
    .B(_02144_),
    .Y(_02235_));
 sky130_fd_sc_hd__mux2_1 _17898_ (.A0(\core.cpuregs[22][20] ),
    .A1(\core.cpuregs[23][20] ),
    .S(_02146_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _17899_ (.A0(\core.cpuregs[20][20] ),
    .A1(\core.cpuregs[21][20] ),
    .S(_02148_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _17900_ (.A0(_02236_),
    .A1(_02237_),
    .S(_02150_),
    .X(_02238_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17901_ (.A(_10369_),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_1 _17902_ (.A(_02238_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__clkbuf_2 _17903_ (.A(_10357_),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _17904_ (.A0(\core.cpuregs[6][20] ),
    .A1(\core.cpuregs[7][20] ),
    .S(_02058_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _17905_ (.A0(\core.cpuregs[4][20] ),
    .A1(\core.cpuregs[5][20] ),
    .S(_02060_),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _17906_ (.A0(_02242_),
    .A1(_02243_),
    .S(_02155_),
    .X(_02244_));
 sky130_fd_sc_hd__clkbuf_4 _17907_ (.A(_09648_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_2 _17908_ (.A0(\core.cpuregs[0][20] ),
    .A1(\core.cpuregs[1][20] ),
    .S(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_4 _17909_ (.A(_10338_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _17910_ (.A0(\core.cpuregs[2][20] ),
    .A1(\core.cpuregs[3][20] ),
    .S(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _17911_ (.A0(_02246_),
    .A1(_02248_),
    .S(_02108_),
    .X(_02249_));
 sky130_fd_sc_hd__buf_1 _17912_ (.A(_04550_),
    .X(_02250_));
 sky130_fd_sc_hd__and2_1 _17913_ (.A(_02249_),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__a211oi_1 _17914_ (.A1(_02241_),
    .A2(_02244_),
    .B1(_02157_),
    .C1(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__a31o_1 _17915_ (.A1(_02094_),
    .A2(_02235_),
    .A3(_02240_),
    .B1(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__nand2_1 _17916_ (.A(_02253_),
    .B(_02022_),
    .Y(_02254_));
 sky130_fd_sc_hd__a22o_1 _17917_ (.A1(\core.decoded_imm[20] ),
    .A2(_02168_),
    .B1(_02231_),
    .B2(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _17918_ (.A0(_02255_),
    .A1(\core.pcpi_rs2[20] ),
    .S(_02166_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _17919_ (.A(_02256_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _17920_ (.A0(\core.cpuregs[24][21] ),
    .A1(\core.cpuregs[25][21] ),
    .S(_02026_),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _17921_ (.A0(\core.cpuregs[26][21] ),
    .A1(\core.cpuregs[27][21] ),
    .S(_02028_),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_2 _17922_ (.A(_04641_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(_02257_),
    .A1(_02258_),
    .S(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_02260_),
    .B(_02076_),
    .Y(_02261_));
 sky130_fd_sc_hd__mux2_1 _17925_ (.A0(\core.cpuregs[28][21] ),
    .A1(\core.cpuregs[29][21] ),
    .S(_02032_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _17926_ (.A0(\core.cpuregs[30][21] ),
    .A1(\core.cpuregs[31][21] ),
    .S(_02034_),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _17927_ (.A0(_02262_),
    .A1(_02263_),
    .S(_02122_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _17928_ (.A(_02264_),
    .B(_02217_),
    .Y(_02265_));
 sky130_fd_sc_hd__mux2_1 _17929_ (.A0(\core.cpuregs[12][21] ),
    .A1(\core.cpuregs[13][21] ),
    .S(_02219_),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _17930_ (.A0(\core.cpuregs[14][21] ),
    .A1(\core.cpuregs[15][21] ),
    .S(_02178_),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _17931_ (.A0(_02266_),
    .A1(_02267_),
    .S(_02084_),
    .X(_02268_));
 sky130_fd_sc_hd__nand2_1 _17932_ (.A(_02268_),
    .B(_02181_),
    .Y(_02269_));
 sky130_fd_sc_hd__mux2_1 _17933_ (.A0(\core.cpuregs[8][21] ),
    .A1(\core.cpuregs[9][21] ),
    .S(_02129_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _17934_ (.A0(\core.cpuregs[10][21] ),
    .A1(\core.cpuregs[11][21] ),
    .S(_02131_),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _17935_ (.A0(_02270_),
    .A1(_02271_),
    .S(_02044_),
    .X(_02272_));
 sky130_fd_sc_hd__nand2_1 _17936_ (.A(_02272_),
    .B(_02227_),
    .Y(_02273_));
 sky130_fd_sc_hd__and3_1 _17937_ (.A(_02269_),
    .B(_02273_),
    .C(_02135_),
    .X(_02274_));
 sky130_fd_sc_hd__a31o_1 _17938_ (.A1(_02072_),
    .A2(_02261_),
    .A3(_02265_),
    .B1(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__clkbuf_4 _17939_ (.A(_04552_),
    .X(_02276_));
 sky130_fd_sc_hd__buf_2 _17940_ (.A(_10385_),
    .X(_02277_));
 sky130_fd_sc_hd__a21oi_4 _17941_ (.A1(_02275_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(\core.cpuregs[16][21] ),
    .A1(\core.cpuregs[17][21] ),
    .S(_02139_),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _17943_ (.A0(\core.cpuregs[18][21] ),
    .A1(\core.cpuregs[19][21] ),
    .S(_02141_),
    .X(_02280_));
 sky130_fd_sc_hd__clkbuf_2 _17944_ (.A(_10395_),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_2 _17945_ (.A0(_02279_),
    .A1(_02280_),
    .S(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__nand2_2 _17946_ (.A(_02282_),
    .B(_02144_),
    .Y(_02283_));
 sky130_fd_sc_hd__mux2_1 _17947_ (.A0(\core.cpuregs[22][21] ),
    .A1(\core.cpuregs[23][21] ),
    .S(_02146_),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _17948_ (.A0(\core.cpuregs[20][21] ),
    .A1(\core.cpuregs[21][21] ),
    .S(_02148_),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _17949_ (.A0(_02284_),
    .A1(_02285_),
    .S(_02150_),
    .X(_02286_));
 sky130_fd_sc_hd__nand2_1 _17950_ (.A(_02286_),
    .B(_02239_),
    .Y(_02287_));
 sky130_fd_sc_hd__mux2_1 _17951_ (.A0(\core.cpuregs[6][21] ),
    .A1(\core.cpuregs[7][21] ),
    .S(_02058_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _17952_ (.A0(\core.cpuregs[4][21] ),
    .A1(\core.cpuregs[5][21] ),
    .S(_02060_),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_2 _17953_ (.A0(_02288_),
    .A1(_02289_),
    .S(_02155_),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _17954_ (.A0(\core.cpuregs[0][21] ),
    .A1(\core.cpuregs[1][21] ),
    .S(_02245_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _17955_ (.A0(\core.cpuregs[2][21] ),
    .A1(\core.cpuregs[3][21] ),
    .S(_02247_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _17956_ (.A0(_02291_),
    .A1(_02292_),
    .S(_02108_),
    .X(_02293_));
 sky130_fd_sc_hd__and2_1 _17957_ (.A(_02293_),
    .B(_02250_),
    .X(_02294_));
 sky130_fd_sc_hd__a211oi_2 _17958_ (.A1(_02241_),
    .A2(_02290_),
    .B1(_02157_),
    .C1(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__a31o_1 _17959_ (.A1(_02094_),
    .A2(_02283_),
    .A3(_02287_),
    .B1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _17960_ (.A(_01746_),
    .X(_02297_));
 sky130_fd_sc_hd__nand2_1 _17961_ (.A(_02296_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__a22o_1 _17962_ (.A1(\core.decoded_imm[21] ),
    .A2(_02168_),
    .B1(_02278_),
    .B2(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _17963_ (.A0(_02299_),
    .A1(\core.pcpi_rs2[21] ),
    .S(_02166_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_1 _17964_ (.A(_02300_),
    .X(_00625_));
 sky130_fd_sc_hd__clkbuf_2 _17965_ (.A(_04567_),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_2 _17966_ (.A0(\core.cpuregs[24][22] ),
    .A1(\core.cpuregs[25][22] ),
    .S(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__clkbuf_2 _17967_ (.A(_04636_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _17968_ (.A0(\core.cpuregs[26][22] ),
    .A1(\core.cpuregs[27][22] ),
    .S(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _17969_ (.A0(_02302_),
    .A1(_02304_),
    .S(_02259_),
    .X(_02305_));
 sky130_fd_sc_hd__nand2_2 _17970_ (.A(_02305_),
    .B(_02076_),
    .Y(_02306_));
 sky130_fd_sc_hd__clkbuf_2 _17971_ (.A(_04662_),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_1 _17972_ (.A0(\core.cpuregs[28][22] ),
    .A1(\core.cpuregs[29][22] ),
    .S(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__buf_4 _17973_ (.A(_10352_),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _17974_ (.A0(\core.cpuregs[30][22] ),
    .A1(\core.cpuregs[31][22] ),
    .S(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _17975_ (.A0(_02308_),
    .A1(_02310_),
    .S(_02122_),
    .X(_02311_));
 sky130_fd_sc_hd__nand2_1 _17976_ (.A(_02311_),
    .B(_02217_),
    .Y(_02312_));
 sky130_fd_sc_hd__mux2_1 _17977_ (.A0(\core.cpuregs[12][22] ),
    .A1(\core.cpuregs[13][22] ),
    .S(_02219_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _17978_ (.A0(\core.cpuregs[14][22] ),
    .A1(\core.cpuregs[15][22] ),
    .S(_02178_),
    .X(_02314_));
 sky130_fd_sc_hd__mux2_1 _17979_ (.A0(_02313_),
    .A1(_02314_),
    .S(_02084_),
    .X(_02315_));
 sky130_fd_sc_hd__nand2_1 _17980_ (.A(_02315_),
    .B(_02181_),
    .Y(_02316_));
 sky130_fd_sc_hd__mux2_1 _17981_ (.A0(\core.cpuregs[8][22] ),
    .A1(\core.cpuregs[9][22] ),
    .S(_02129_),
    .X(_02317_));
 sky130_fd_sc_hd__mux2_1 _17982_ (.A0(\core.cpuregs[10][22] ),
    .A1(\core.cpuregs[11][22] ),
    .S(_02131_),
    .X(_02318_));
 sky130_fd_sc_hd__clkbuf_4 _17983_ (.A(_04640_),
    .X(_02319_));
 sky130_fd_sc_hd__mux2_1 _17984_ (.A0(_02317_),
    .A1(_02318_),
    .S(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(_02320_),
    .B(_02227_),
    .Y(_02321_));
 sky130_fd_sc_hd__and3_1 _17986_ (.A(_02316_),
    .B(_02321_),
    .C(_02135_),
    .X(_02322_));
 sky130_fd_sc_hd__a31o_1 _17987_ (.A1(_02072_),
    .A2(_02306_),
    .A3(_02312_),
    .B1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__a21oi_1 _17988_ (.A1(_02323_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02324_));
 sky130_fd_sc_hd__mux2_1 _17989_ (.A0(\core.cpuregs[16][22] ),
    .A1(\core.cpuregs[17][22] ),
    .S(_02139_),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _17990_ (.A0(\core.cpuregs[18][22] ),
    .A1(\core.cpuregs[19][22] ),
    .S(_02141_),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _17991_ (.A0(_02325_),
    .A1(_02326_),
    .S(_02281_),
    .X(_02327_));
 sky130_fd_sc_hd__nand2_2 _17992_ (.A(_02327_),
    .B(_02144_),
    .Y(_02328_));
 sky130_fd_sc_hd__mux2_1 _17993_ (.A0(\core.cpuregs[22][22] ),
    .A1(\core.cpuregs[23][22] ),
    .S(_02146_),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _17994_ (.A0(\core.cpuregs[20][22] ),
    .A1(\core.cpuregs[21][22] ),
    .S(_02148_),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _17995_ (.A0(_02329_),
    .A1(_02330_),
    .S(_02150_),
    .X(_02331_));
 sky130_fd_sc_hd__nand2_1 _17996_ (.A(_02331_),
    .B(_02239_),
    .Y(_02332_));
 sky130_fd_sc_hd__clkbuf_4 _17997_ (.A(_10413_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _17998_ (.A0(\core.cpuregs[6][22] ),
    .A1(\core.cpuregs[7][22] ),
    .S(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__clkbuf_4 _17999_ (.A(_10413_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _18000_ (.A0(\core.cpuregs[4][22] ),
    .A1(\core.cpuregs[5][22] ),
    .S(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _18001_ (.A0(_02334_),
    .A1(_02336_),
    .S(_02155_),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _18002_ (.A0(\core.cpuregs[0][22] ),
    .A1(\core.cpuregs[1][22] ),
    .S(_02245_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _18003_ (.A0(\core.cpuregs[2][22] ),
    .A1(\core.cpuregs[3][22] ),
    .S(_02247_),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _18004_ (.A0(_02338_),
    .A1(_02339_),
    .S(_02108_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_1 _18005_ (.A(_02340_),
    .B(_02250_),
    .X(_02341_));
 sky130_fd_sc_hd__a211oi_1 _18006_ (.A1(_02241_),
    .A2(_02337_),
    .B1(_02157_),
    .C1(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__a31o_1 _18007_ (.A1(_02094_),
    .A2(_02328_),
    .A3(_02332_),
    .B1(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__nand2_1 _18008_ (.A(_02343_),
    .B(_02297_),
    .Y(_02344_));
 sky130_fd_sc_hd__a22o_1 _18009_ (.A1(\core.decoded_imm[22] ),
    .A2(_02168_),
    .B1(_02324_),
    .B2(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_2 _18010_ (.A0(_02345_),
    .A1(\core.pcpi_rs2[22] ),
    .S(_02166_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_2 _18011_ (.A(_02346_),
    .X(_00626_));
 sky130_fd_sc_hd__clkbuf_4 _18012_ (.A(_10418_),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_4 _18013_ (.A0(\core.cpuregs[24][23] ),
    .A1(\core.cpuregs[25][23] ),
    .S(_02301_),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_4 _18014_ (.A0(\core.cpuregs[26][23] ),
    .A1(\core.cpuregs[27][23] ),
    .S(_02303_),
    .X(_02349_));
 sky130_fd_sc_hd__mux2_1 _18015_ (.A0(_02348_),
    .A1(_02349_),
    .S(_02259_),
    .X(_02350_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18016_ (.A(_10347_),
    .X(_02351_));
 sky130_fd_sc_hd__nand2_1 _18017_ (.A(_02350_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__mux2_1 _18018_ (.A0(\core.cpuregs[28][23] ),
    .A1(\core.cpuregs[29][23] ),
    .S(_02307_),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_4 _18019_ (.A0(\core.cpuregs[30][23] ),
    .A1(\core.cpuregs[31][23] ),
    .S(_02309_),
    .X(_02354_));
 sky130_fd_sc_hd__mux2_1 _18020_ (.A0(_02353_),
    .A1(_02354_),
    .S(_02122_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_1 _18021_ (.A(_02355_),
    .B(_02217_),
    .Y(_02356_));
 sky130_fd_sc_hd__mux2_1 _18022_ (.A0(\core.cpuregs[12][23] ),
    .A1(\core.cpuregs[13][23] ),
    .S(_02219_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _18023_ (.A0(\core.cpuregs[14][23] ),
    .A1(\core.cpuregs[15][23] ),
    .S(_02178_),
    .X(_02358_));
 sky130_fd_sc_hd__clkbuf_4 _18024_ (.A(_10365_),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_4 _18025_ (.A0(_02357_),
    .A1(_02358_),
    .S(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(_02360_),
    .B(_02181_),
    .Y(_02361_));
 sky130_fd_sc_hd__mux2_1 _18027_ (.A0(\core.cpuregs[8][23] ),
    .A1(\core.cpuregs[9][23] ),
    .S(_02129_),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _18028_ (.A0(\core.cpuregs[10][23] ),
    .A1(\core.cpuregs[11][23] ),
    .S(_02131_),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _18029_ (.A0(_02362_),
    .A1(_02363_),
    .S(_02319_),
    .X(_02364_));
 sky130_fd_sc_hd__nand2_1 _18030_ (.A(_02364_),
    .B(_02227_),
    .Y(_02365_));
 sky130_fd_sc_hd__and3_1 _18031_ (.A(_02361_),
    .B(_02365_),
    .C(_02135_),
    .X(_02366_));
 sky130_fd_sc_hd__a31o_1 _18032_ (.A1(_02347_),
    .A2(_02352_),
    .A3(_02356_),
    .B1(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a21oi_4 _18033_ (.A1(_02367_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02368_));
 sky130_fd_sc_hd__clkbuf_4 _18034_ (.A(_10336_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _18035_ (.A0(\core.cpuregs[16][23] ),
    .A1(\core.cpuregs[17][23] ),
    .S(_02139_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _18036_ (.A0(\core.cpuregs[18][23] ),
    .A1(\core.cpuregs[19][23] ),
    .S(_02141_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _18037_ (.A0(_02370_),
    .A1(_02371_),
    .S(_02281_),
    .X(_02372_));
 sky130_fd_sc_hd__nand2_1 _18038_ (.A(_02372_),
    .B(_02144_),
    .Y(_02373_));
 sky130_fd_sc_hd__mux2_1 _18039_ (.A0(\core.cpuregs[22][23] ),
    .A1(\core.cpuregs[23][23] ),
    .S(_02146_),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_2 _18040_ (.A0(\core.cpuregs[20][23] ),
    .A1(\core.cpuregs[21][23] ),
    .S(_02148_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _18041_ (.A0(_02374_),
    .A1(_02375_),
    .S(_02150_),
    .X(_02376_));
 sky130_fd_sc_hd__nand2_1 _18042_ (.A(_02376_),
    .B(_02239_),
    .Y(_02377_));
 sky130_fd_sc_hd__mux2_1 _18043_ (.A0(\core.cpuregs[6][23] ),
    .A1(\core.cpuregs[7][23] ),
    .S(_02333_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _18044_ (.A0(\core.cpuregs[4][23] ),
    .A1(\core.cpuregs[5][23] ),
    .S(_02335_),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _18045_ (.A0(_02378_),
    .A1(_02379_),
    .S(_02155_),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _18046_ (.A0(\core.cpuregs[0][23] ),
    .A1(\core.cpuregs[1][23] ),
    .S(_02245_),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _18047_ (.A0(\core.cpuregs[2][23] ),
    .A1(\core.cpuregs[3][23] ),
    .S(_02247_),
    .X(_02382_));
 sky130_fd_sc_hd__clkbuf_2 _18048_ (.A(_10365_),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _18049_ (.A0(_02381_),
    .A1(_02382_),
    .S(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__and2_1 _18050_ (.A(_02384_),
    .B(_02250_),
    .X(_02385_));
 sky130_fd_sc_hd__a211oi_2 _18051_ (.A1(_02241_),
    .A2(_02380_),
    .B1(_02157_),
    .C1(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__a31o_1 _18052_ (.A1(_02369_),
    .A2(_02373_),
    .A3(_02377_),
    .B1(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__nand2_1 _18053_ (.A(_02387_),
    .B(_02297_),
    .Y(_02388_));
 sky130_fd_sc_hd__a22o_1 _18054_ (.A1(\core.decoded_imm[23] ),
    .A2(_02168_),
    .B1(_02368_),
    .B2(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _18055_ (.A0(_02389_),
    .A1(\core.pcpi_rs2[23] ),
    .S(_02166_),
    .X(_02390_));
 sky130_fd_sc_hd__clkbuf_1 _18056_ (.A(_02390_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _18057_ (.A0(\core.cpuregs[24][24] ),
    .A1(\core.cpuregs[25][24] ),
    .S(_02301_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_2 _18058_ (.A0(\core.cpuregs[26][24] ),
    .A1(\core.cpuregs[27][24] ),
    .S(_02303_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_2 _18059_ (.A0(_02391_),
    .A1(_02392_),
    .S(_02259_),
    .X(_02393_));
 sky130_fd_sc_hd__nand2_1 _18060_ (.A(_02393_),
    .B(_02351_),
    .Y(_02394_));
 sky130_fd_sc_hd__mux2_1 _18061_ (.A0(\core.cpuregs[28][24] ),
    .A1(\core.cpuregs[29][24] ),
    .S(_02307_),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_2 _18062_ (.A0(\core.cpuregs[30][24] ),
    .A1(\core.cpuregs[31][24] ),
    .S(_02309_),
    .X(_02396_));
 sky130_fd_sc_hd__clkbuf_2 _18063_ (.A(_09617_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _18064_ (.A0(_02395_),
    .A1(_02396_),
    .S(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(_02398_),
    .B(_02217_),
    .Y(_02399_));
 sky130_fd_sc_hd__mux2_1 _18066_ (.A0(\core.cpuregs[12][24] ),
    .A1(\core.cpuregs[13][24] ),
    .S(_02219_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _18067_ (.A0(\core.cpuregs[14][24] ),
    .A1(\core.cpuregs[15][24] ),
    .S(_02178_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_2 _18068_ (.A0(_02400_),
    .A1(_02401_),
    .S(_02359_),
    .X(_02402_));
 sky130_fd_sc_hd__nand2_1 _18069_ (.A(_02402_),
    .B(_02181_),
    .Y(_02403_));
 sky130_fd_sc_hd__clkbuf_4 _18070_ (.A(_04521_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_4 _18071_ (.A0(\core.cpuregs[8][24] ),
    .A1(\core.cpuregs[9][24] ),
    .S(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__clkbuf_2 _18072_ (.A(_04521_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _18073_ (.A0(\core.cpuregs[10][24] ),
    .A1(\core.cpuregs[11][24] ),
    .S(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _18074_ (.A0(_02405_),
    .A1(_02407_),
    .S(_02319_),
    .X(_02408_));
 sky130_fd_sc_hd__nand2_1 _18075_ (.A(_02408_),
    .B(_02227_),
    .Y(_02409_));
 sky130_fd_sc_hd__buf_2 _18076_ (.A(_10379_),
    .X(_02410_));
 sky130_fd_sc_hd__and3_1 _18077_ (.A(_02403_),
    .B(_02409_),
    .C(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__a31o_1 _18078_ (.A1(_02347_),
    .A2(_02394_),
    .A3(_02399_),
    .B1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a21oi_1 _18079_ (.A1(_02412_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02413_));
 sky130_fd_sc_hd__clkbuf_2 _18080_ (.A(_10339_),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _18081_ (.A0(\core.cpuregs[16][24] ),
    .A1(\core.cpuregs[17][24] ),
    .S(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__clkbuf_2 _18082_ (.A(_10392_),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _18083_ (.A0(\core.cpuregs[18][24] ),
    .A1(\core.cpuregs[19][24] ),
    .S(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _18084_ (.A0(_02415_),
    .A1(_02417_),
    .S(_02281_),
    .X(_02418_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18085_ (.A(_10399_),
    .X(_02419_));
 sky130_fd_sc_hd__nand2_1 _18086_ (.A(_02418_),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__clkbuf_2 _18087_ (.A(_04522_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _18088_ (.A0(\core.cpuregs[22][24] ),
    .A1(\core.cpuregs[23][24] ),
    .S(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__buf_4 _18089_ (.A(_04532_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _18090_ (.A0(\core.cpuregs[20][24] ),
    .A1(\core.cpuregs[21][24] ),
    .S(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__clkbuf_2 _18091_ (.A(_04537_),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _18092_ (.A0(_02422_),
    .A1(_02424_),
    .S(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_1 _18093_ (.A(_02426_),
    .B(_02239_),
    .Y(_02427_));
 sky130_fd_sc_hd__mux2_2 _18094_ (.A0(\core.cpuregs[6][24] ),
    .A1(\core.cpuregs[7][24] ),
    .S(_02333_),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _18095_ (.A0(\core.cpuregs[4][24] ),
    .A1(\core.cpuregs[5][24] ),
    .S(_02335_),
    .X(_02429_));
 sky130_fd_sc_hd__clkbuf_4 _18096_ (.A(_09622_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _18097_ (.A0(_02428_),
    .A1(_02429_),
    .S(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_2 _18098_ (.A(_00004_),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _18099_ (.A0(\core.cpuregs[0][24] ),
    .A1(\core.cpuregs[1][24] ),
    .S(_02245_),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_2 _18100_ (.A0(\core.cpuregs[2][24] ),
    .A1(\core.cpuregs[3][24] ),
    .S(_02247_),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _18101_ (.A0(_02433_),
    .A1(_02434_),
    .S(_02383_),
    .X(_02435_));
 sky130_fd_sc_hd__and2_1 _18102_ (.A(_02435_),
    .B(_02250_),
    .X(_02436_));
 sky130_fd_sc_hd__a211oi_1 _18103_ (.A1(_02241_),
    .A2(_02431_),
    .B1(_02432_),
    .C1(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a31o_1 _18104_ (.A1(_02369_),
    .A2(_02420_),
    .A3(_02427_),
    .B1(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_1 _18105_ (.A(_02438_),
    .B(_02297_),
    .Y(_02439_));
 sky130_fd_sc_hd__a22o_1 _18106_ (.A1(\core.decoded_imm[24] ),
    .A2(_02168_),
    .B1(_02413_),
    .B2(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__clkbuf_4 _18107_ (.A(_10321_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _18108_ (.A0(_02440_),
    .A1(\core.pcpi_rs2[24] ),
    .S(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__clkbuf_1 _18109_ (.A(_02442_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _18110_ (.A0(\core.cpuregs[24][25] ),
    .A1(\core.cpuregs[25][25] ),
    .S(_02301_),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _18111_ (.A0(\core.cpuregs[26][25] ),
    .A1(\core.cpuregs[27][25] ),
    .S(_02303_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_2 _18112_ (.A0(_02443_),
    .A1(_02444_),
    .S(_02259_),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_1 _18113_ (.A(_02445_),
    .B(_02351_),
    .Y(_02446_));
 sky130_fd_sc_hd__mux2_1 _18114_ (.A0(\core.cpuregs[28][25] ),
    .A1(\core.cpuregs[29][25] ),
    .S(_02307_),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _18115_ (.A0(\core.cpuregs[30][25] ),
    .A1(\core.cpuregs[31][25] ),
    .S(_02309_),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _18116_ (.A0(_02447_),
    .A1(_02448_),
    .S(_02397_),
    .X(_02449_));
 sky130_fd_sc_hd__nand2_1 _18117_ (.A(_02449_),
    .B(_02217_),
    .Y(_02450_));
 sky130_fd_sc_hd__mux2_1 _18118_ (.A0(\core.cpuregs[12][25] ),
    .A1(\core.cpuregs[13][25] ),
    .S(_02219_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _18119_ (.A0(\core.cpuregs[14][25] ),
    .A1(\core.cpuregs[15][25] ),
    .S(_01670_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _18120_ (.A0(_02451_),
    .A1(_02452_),
    .S(_02359_),
    .X(_02453_));
 sky130_fd_sc_hd__nand2_1 _18121_ (.A(_02453_),
    .B(_01632_),
    .Y(_02454_));
 sky130_fd_sc_hd__mux2_1 _18122_ (.A0(\core.cpuregs[8][25] ),
    .A1(\core.cpuregs[9][25] ),
    .S(_02404_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _18123_ (.A0(\core.cpuregs[10][25] ),
    .A1(\core.cpuregs[11][25] ),
    .S(_02406_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _18124_ (.A0(_02455_),
    .A1(_02456_),
    .S(_02319_),
    .X(_02457_));
 sky130_fd_sc_hd__nand2_1 _18125_ (.A(_02457_),
    .B(_02227_),
    .Y(_02458_));
 sky130_fd_sc_hd__and3_1 _18126_ (.A(_02454_),
    .B(_02458_),
    .C(_02410_),
    .X(_02459_));
 sky130_fd_sc_hd__a31o_1 _18127_ (.A1(_02347_),
    .A2(_02446_),
    .A3(_02450_),
    .B1(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__a21oi_1 _18128_ (.A1(_02460_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02461_));
 sky130_fd_sc_hd__mux2_1 _18129_ (.A0(\core.cpuregs[16][25] ),
    .A1(\core.cpuregs[17][25] ),
    .S(_02414_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _18130_ (.A0(\core.cpuregs[18][25] ),
    .A1(\core.cpuregs[19][25] ),
    .S(_02416_),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _18131_ (.A0(_02462_),
    .A1(_02463_),
    .S(_02281_),
    .X(_02464_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(_02464_),
    .B(_02419_),
    .Y(_02465_));
 sky130_fd_sc_hd__mux2_1 _18133_ (.A0(\core.cpuregs[22][25] ),
    .A1(\core.cpuregs[23][25] ),
    .S(_02421_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _18134_ (.A0(\core.cpuregs[20][25] ),
    .A1(\core.cpuregs[21][25] ),
    .S(_02423_),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _18135_ (.A0(_02466_),
    .A1(_02467_),
    .S(_02425_),
    .X(_02468_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_02468_),
    .B(_02239_),
    .Y(_02469_));
 sky130_fd_sc_hd__mux2_1 _18137_ (.A0(\core.cpuregs[6][25] ),
    .A1(\core.cpuregs[7][25] ),
    .S(_02333_),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _18138_ (.A0(\core.cpuregs[4][25] ),
    .A1(\core.cpuregs[5][25] ),
    .S(_02335_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _18139_ (.A0(_02470_),
    .A1(_02471_),
    .S(_02430_),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _18140_ (.A0(\core.cpuregs[0][25] ),
    .A1(\core.cpuregs[1][25] ),
    .S(_02245_),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _18141_ (.A0(\core.cpuregs[2][25] ),
    .A1(\core.cpuregs[3][25] ),
    .S(_02247_),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_2 _18142_ (.A0(_02473_),
    .A1(_02474_),
    .S(_02383_),
    .X(_02475_));
 sky130_fd_sc_hd__and2_1 _18143_ (.A(_02475_),
    .B(_02250_),
    .X(_02476_));
 sky130_fd_sc_hd__a211oi_1 _18144_ (.A1(_02241_),
    .A2(_02472_),
    .B1(_02432_),
    .C1(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a31o_1 _18145_ (.A1(_02369_),
    .A2(_02465_),
    .A3(_02469_),
    .B1(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__nand2_1 _18146_ (.A(_02478_),
    .B(_02297_),
    .Y(_02479_));
 sky130_fd_sc_hd__a22o_1 _18147_ (.A1(\core.decoded_imm[25] ),
    .A2(_04497_),
    .B1(_02461_),
    .B2(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _18148_ (.A0(_02480_),
    .A1(\core.pcpi_rs2[25] ),
    .S(_02441_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_1 _18149_ (.A(_02481_),
    .X(_00629_));
 sky130_fd_sc_hd__o21ai_2 _18150_ (.A1(_06190_),
    .A2(_04474_),
    .B1(_01649_),
    .Y(_02482_));
 sky130_fd_sc_hd__mux2_1 _18151_ (.A0(\core.cpuregs[16][26] ),
    .A1(\core.cpuregs[17][26] ),
    .S(_01652_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_2 _18152_ (.A0(\core.cpuregs[18][26] ),
    .A1(\core.cpuregs[19][26] ),
    .S(_01652_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _18153_ (.A0(_02483_),
    .A1(_02484_),
    .S(_01655_),
    .X(_02485_));
 sky130_fd_sc_hd__nand2_1 _18154_ (.A(_02485_),
    .B(_01657_),
    .Y(_02486_));
 sky130_fd_sc_hd__mux2_1 _18155_ (.A0(\core.cpuregs[22][26] ),
    .A1(\core.cpuregs[23][26] ),
    .S(_01659_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _18156_ (.A0(\core.cpuregs[20][26] ),
    .A1(\core.cpuregs[21][26] ),
    .S(_01659_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _18157_ (.A0(_02487_),
    .A1(_02488_),
    .S(_01662_),
    .X(_02489_));
 sky130_fd_sc_hd__nand2_1 _18158_ (.A(_02489_),
    .B(_01664_),
    .Y(_02490_));
 sky130_fd_sc_hd__mux2_1 _18159_ (.A0(\core.cpuregs[6][26] ),
    .A1(\core.cpuregs[7][26] ),
    .S(_01666_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _18160_ (.A0(\core.cpuregs[4][26] ),
    .A1(\core.cpuregs[5][26] ),
    .S(_01666_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _18161_ (.A0(_02491_),
    .A1(_02492_),
    .S(_01662_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _18162_ (.A0(\core.cpuregs[0][26] ),
    .A1(\core.cpuregs[1][26] ),
    .S(_01671_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _18163_ (.A0(\core.cpuregs[2][26] ),
    .A1(\core.cpuregs[3][26] ),
    .S(_01671_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _18164_ (.A0(_02494_),
    .A1(_02495_),
    .S(_01674_),
    .X(_02496_));
 sky130_fd_sc_hd__and2_1 _18165_ (.A(_02496_),
    .B(_01676_),
    .X(_02497_));
 sky130_fd_sc_hd__a211oi_1 _18166_ (.A1(_01664_),
    .A2(_02493_),
    .B1(_01651_),
    .C1(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__a31o_1 _18167_ (.A1(_01651_),
    .A2(_02486_),
    .A3(_02490_),
    .B1(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _18168_ (.A0(\core.cpuregs[24][26] ),
    .A1(\core.cpuregs[25][26] ),
    .S(_01681_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _18169_ (.A0(\core.cpuregs[26][26] ),
    .A1(\core.cpuregs[27][26] ),
    .S(_01681_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_8 _18170_ (.A0(_02500_),
    .A1(_02501_),
    .S(_01655_),
    .X(_02502_));
 sky130_fd_sc_hd__nand2_1 _18171_ (.A(_02502_),
    .B(_01657_),
    .Y(_02503_));
 sky130_fd_sc_hd__mux2_1 _18172_ (.A0(\core.cpuregs[28][26] ),
    .A1(\core.cpuregs[29][26] ),
    .S(_01686_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _18173_ (.A0(\core.cpuregs[30][26] ),
    .A1(\core.cpuregs[31][26] ),
    .S(_01686_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_8 _18174_ (.A0(_02504_),
    .A1(_02505_),
    .S(_01674_),
    .X(_02506_));
 sky130_fd_sc_hd__nand2_1 _18175_ (.A(_02506_),
    .B(_10408_),
    .Y(_02507_));
 sky130_fd_sc_hd__mux2_1 _18176_ (.A0(\core.cpuregs[8][26] ),
    .A1(\core.cpuregs[9][26] ),
    .S(_01691_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _18177_ (.A0(\core.cpuregs[10][26] ),
    .A1(\core.cpuregs[11][26] ),
    .S(_01691_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _18178_ (.A0(_02508_),
    .A1(_02509_),
    .S(_10396_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _18179_ (.A0(\core.cpuregs[12][26] ),
    .A1(\core.cpuregs[13][26] ),
    .S(_01695_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _18180_ (.A0(\core.cpuregs[14][26] ),
    .A1(\core.cpuregs[15][26] ),
    .S(_10350_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _18181_ (.A0(_02511_),
    .A1(_02512_),
    .S(_01698_),
    .X(_02513_));
 sky130_fd_sc_hd__and2_1 _18182_ (.A(_02513_),
    .B(_01700_),
    .X(_02514_));
 sky130_fd_sc_hd__a211oi_1 _18183_ (.A1(_01676_),
    .A2(_02510_),
    .B1(_01680_),
    .C1(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__a31o_1 _18184_ (.A1(_01680_),
    .A2(_02503_),
    .A3(_02507_),
    .B1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_1 _18185_ (.A1(_02516_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_02517_));
 sky130_fd_sc_hd__a21boi_1 _18186_ (.A1(_10431_),
    .A2(_02499_),
    .B1_N(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__o22a_1 _18187_ (.A1(\core.pcpi_rs2[26] ),
    .A2(_01649_),
    .B1(_02482_),
    .B2(_02518_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _18188_ (.A0(\core.cpuregs[24][27] ),
    .A1(\core.cpuregs[25][27] ),
    .S(_02301_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _18189_ (.A0(\core.cpuregs[26][27] ),
    .A1(\core.cpuregs[27][27] ),
    .S(_02303_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_2 _18190_ (.A0(_02519_),
    .A1(_02520_),
    .S(_02259_),
    .X(_02521_));
 sky130_fd_sc_hd__nand2_1 _18191_ (.A(_02521_),
    .B(_02351_),
    .Y(_02522_));
 sky130_fd_sc_hd__mux2_2 _18192_ (.A0(\core.cpuregs[28][27] ),
    .A1(\core.cpuregs[29][27] ),
    .S(_02307_),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _18193_ (.A0(\core.cpuregs[30][27] ),
    .A1(\core.cpuregs[31][27] ),
    .S(_02309_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _18194_ (.A0(_02523_),
    .A1(_02524_),
    .S(_02397_),
    .X(_02525_));
 sky130_fd_sc_hd__nand2_1 _18195_ (.A(_02525_),
    .B(_01700_),
    .Y(_02526_));
 sky130_fd_sc_hd__mux2_1 _18196_ (.A0(\core.cpuregs[12][27] ),
    .A1(\core.cpuregs[13][27] ),
    .S(_10363_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _18197_ (.A0(\core.cpuregs[14][27] ),
    .A1(\core.cpuregs[15][27] ),
    .S(_01670_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _18198_ (.A0(_02527_),
    .A1(_02528_),
    .S(_02359_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _18199_ (.A(_02529_),
    .B(_01632_),
    .Y(_02530_));
 sky130_fd_sc_hd__mux2_1 _18200_ (.A0(\core.cpuregs[8][27] ),
    .A1(\core.cpuregs[9][27] ),
    .S(_02404_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_4 _18201_ (.A0(\core.cpuregs[10][27] ),
    .A1(\core.cpuregs[11][27] ),
    .S(_02406_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _18202_ (.A0(_02531_),
    .A1(_02532_),
    .S(_02319_),
    .X(_02533_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(_02533_),
    .B(_10426_),
    .Y(_02534_));
 sky130_fd_sc_hd__and3_1 _18204_ (.A(_02530_),
    .B(_02534_),
    .C(_02410_),
    .X(_02535_));
 sky130_fd_sc_hd__a31o_1 _18205_ (.A1(_02347_),
    .A2(_02522_),
    .A3(_02526_),
    .B1(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__a21oi_1 _18206_ (.A1(_02536_),
    .A2(_02276_),
    .B1(_02277_),
    .Y(_02537_));
 sky130_fd_sc_hd__mux2_1 _18207_ (.A0(\core.cpuregs[16][27] ),
    .A1(\core.cpuregs[17][27] ),
    .S(_02414_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _18208_ (.A0(\core.cpuregs[18][27] ),
    .A1(\core.cpuregs[19][27] ),
    .S(_02416_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _18209_ (.A0(_02538_),
    .A1(_02539_),
    .S(_02281_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _18210_ (.A(_02540_),
    .B(_02419_),
    .Y(_02541_));
 sky130_fd_sc_hd__mux2_1 _18211_ (.A0(\core.cpuregs[22][27] ),
    .A1(\core.cpuregs[23][27] ),
    .S(_02421_),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _18212_ (.A0(\core.cpuregs[20][27] ),
    .A1(\core.cpuregs[21][27] ),
    .S(_02423_),
    .X(_02543_));
 sky130_fd_sc_hd__mux2_1 _18213_ (.A0(_02542_),
    .A1(_02543_),
    .S(_02425_),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_1 _18214_ (.A(_02544_),
    .B(_10410_),
    .Y(_02545_));
 sky130_fd_sc_hd__mux2_1 _18215_ (.A0(\core.cpuregs[6][27] ),
    .A1(\core.cpuregs[7][27] ),
    .S(_02333_),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_1 _18216_ (.A0(\core.cpuregs[4][27] ),
    .A1(\core.cpuregs[5][27] ),
    .S(_02335_),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_2 _18217_ (.A0(_02546_),
    .A1(_02547_),
    .S(_02430_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _18218_ (.A0(\core.cpuregs[0][27] ),
    .A1(\core.cpuregs[1][27] ),
    .S(_10422_),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _18219_ (.A0(\core.cpuregs[2][27] ),
    .A1(\core.cpuregs[3][27] ),
    .S(_10360_),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _18220_ (.A0(_02549_),
    .A1(_02550_),
    .S(_02383_),
    .X(_02551_));
 sky130_fd_sc_hd__and2_1 _18221_ (.A(_02551_),
    .B(_10398_),
    .X(_02552_));
 sky130_fd_sc_hd__a211oi_1 _18222_ (.A1(_10358_),
    .A2(_02548_),
    .B1(_02432_),
    .C1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__a31o_1 _18223_ (.A1(_02369_),
    .A2(_02541_),
    .A3(_02545_),
    .B1(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(_02554_),
    .B(_02297_),
    .Y(_02555_));
 sky130_fd_sc_hd__a22o_1 _18225_ (.A1(\core.decoded_imm[27] ),
    .A2(_04497_),
    .B1(_02537_),
    .B2(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _18226_ (.A0(_02556_),
    .A1(\core.pcpi_rs2[27] ),
    .S(_02441_),
    .X(_02557_));
 sky130_fd_sc_hd__clkbuf_1 _18227_ (.A(_02557_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _18228_ (.A0(\core.cpuregs[24][28] ),
    .A1(\core.cpuregs[25][28] ),
    .S(_02301_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _18229_ (.A0(\core.cpuregs[26][28] ),
    .A1(\core.cpuregs[27][28] ),
    .S(_02303_),
    .X(_02559_));
 sky130_fd_sc_hd__mux2_1 _18230_ (.A0(_02558_),
    .A1(_02559_),
    .S(_01698_),
    .X(_02560_));
 sky130_fd_sc_hd__nand2_1 _18231_ (.A(_02560_),
    .B(_02351_),
    .Y(_02561_));
 sky130_fd_sc_hd__mux2_2 _18232_ (.A0(\core.cpuregs[28][28] ),
    .A1(\core.cpuregs[29][28] ),
    .S(_02307_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_4 _18233_ (.A0(\core.cpuregs[30][28] ),
    .A1(\core.cpuregs[31][28] ),
    .S(_02309_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _18234_ (.A0(_02562_),
    .A1(_02563_),
    .S(_02397_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _18235_ (.A(_02564_),
    .B(_01700_),
    .Y(_02565_));
 sky130_fd_sc_hd__mux2_1 _18236_ (.A0(\core.cpuregs[12][28] ),
    .A1(\core.cpuregs[13][28] ),
    .S(_10363_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _18237_ (.A0(\core.cpuregs[14][28] ),
    .A1(\core.cpuregs[15][28] ),
    .S(_01670_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_2 _18238_ (.A0(_02566_),
    .A1(_02567_),
    .S(_02359_),
    .X(_02568_));
 sky130_fd_sc_hd__nand2_2 _18239_ (.A(_02568_),
    .B(_01632_),
    .Y(_02569_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(\core.cpuregs[8][28] ),
    .A1(\core.cpuregs[9][28] ),
    .S(_02404_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _18241_ (.A0(\core.cpuregs[10][28] ),
    .A1(\core.cpuregs[11][28] ),
    .S(_02406_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _18242_ (.A0(_02570_),
    .A1(_02571_),
    .S(_02319_),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_1 _18243_ (.A(_02572_),
    .B(_10426_),
    .Y(_02573_));
 sky130_fd_sc_hd__and3_1 _18244_ (.A(_02569_),
    .B(_02573_),
    .C(_02410_),
    .X(_02574_));
 sky130_fd_sc_hd__a31o_1 _18245_ (.A1(_02347_),
    .A2(_02561_),
    .A3(_02565_),
    .B1(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__a21oi_4 _18246_ (.A1(_02575_),
    .A2(_10383_),
    .B1(_10386_),
    .Y(_02576_));
 sky130_fd_sc_hd__mux2_1 _18247_ (.A0(\core.cpuregs[16][28] ),
    .A1(\core.cpuregs[17][28] ),
    .S(_02414_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _18248_ (.A0(\core.cpuregs[18][28] ),
    .A1(\core.cpuregs[19][28] ),
    .S(_02416_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_2 _18249_ (.A0(_02577_),
    .A1(_02578_),
    .S(_10344_),
    .X(_02579_));
 sky130_fd_sc_hd__nand2_1 _18250_ (.A(_02579_),
    .B(_02419_),
    .Y(_02580_));
 sky130_fd_sc_hd__mux2_1 _18251_ (.A0(\core.cpuregs[22][28] ),
    .A1(\core.cpuregs[23][28] ),
    .S(_02421_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _18252_ (.A0(\core.cpuregs[20][28] ),
    .A1(\core.cpuregs[21][28] ),
    .S(_02423_),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_2 _18253_ (.A0(_02581_),
    .A1(_02582_),
    .S(_02425_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_2 _18254_ (.A(_02583_),
    .B(_10410_),
    .Y(_02584_));
 sky130_fd_sc_hd__mux2_1 _18255_ (.A0(\core.cpuregs[6][28] ),
    .A1(\core.cpuregs[7][28] ),
    .S(_02333_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _18256_ (.A0(\core.cpuregs[4][28] ),
    .A1(\core.cpuregs[5][28] ),
    .S(_02335_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _18257_ (.A0(_02585_),
    .A1(_02586_),
    .S(_02430_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _18258_ (.A0(\core.cpuregs[0][28] ),
    .A1(\core.cpuregs[1][28] ),
    .S(_10422_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_2 _18259_ (.A0(\core.cpuregs[2][28] ),
    .A1(\core.cpuregs[3][28] ),
    .S(_10360_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _18260_ (.A0(_02588_),
    .A1(_02589_),
    .S(_02383_),
    .X(_02590_));
 sky130_fd_sc_hd__and2_1 _18261_ (.A(_02590_),
    .B(_10398_),
    .X(_02591_));
 sky130_fd_sc_hd__a211oi_2 _18262_ (.A1(_10358_),
    .A2(_02587_),
    .B1(_02432_),
    .C1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__a31o_1 _18263_ (.A1(_02369_),
    .A2(_02580_),
    .A3(_02584_),
    .B1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _18264_ (.A(_02593_),
    .B(_01746_),
    .Y(_02594_));
 sky130_fd_sc_hd__a22o_1 _18265_ (.A1(\core.decoded_imm[28] ),
    .A2(_04497_),
    .B1(_02576_),
    .B2(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _18266_ (.A0(_02595_),
    .A1(\core.pcpi_rs2[28] ),
    .S(_02441_),
    .X(_02596_));
 sky130_fd_sc_hd__clkbuf_1 _18267_ (.A(_02596_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _18268_ (.A0(\core.cpuregs[24][29] ),
    .A1(\core.cpuregs[25][29] ),
    .S(_10342_),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_2 _18269_ (.A0(\core.cpuregs[26][29] ),
    .A1(\core.cpuregs[27][29] ),
    .S(_01695_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _18270_ (.A0(_02597_),
    .A1(_02598_),
    .S(_01698_),
    .X(_02599_));
 sky130_fd_sc_hd__nand2_1 _18271_ (.A(_02599_),
    .B(_02351_),
    .Y(_02600_));
 sky130_fd_sc_hd__mux2_4 _18272_ (.A0(\core.cpuregs[28][29] ),
    .A1(\core.cpuregs[29][29] ),
    .S(_10353_),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_4 _18273_ (.A0(\core.cpuregs[30][29] ),
    .A1(\core.cpuregs[31][29] ),
    .S(_10411_),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_4 _18274_ (.A0(_02601_),
    .A1(_02602_),
    .S(_02397_),
    .X(_02603_));
 sky130_fd_sc_hd__nand2_1 _18275_ (.A(_02603_),
    .B(_01700_),
    .Y(_02604_));
 sky130_fd_sc_hd__mux2_1 _18276_ (.A0(\core.cpuregs[12][29] ),
    .A1(\core.cpuregs[13][29] ),
    .S(_10363_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _18277_ (.A0(\core.cpuregs[14][29] ),
    .A1(\core.cpuregs[15][29] ),
    .S(_01670_),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _18278_ (.A0(_02605_),
    .A1(_02606_),
    .S(_02359_),
    .X(_02607_));
 sky130_fd_sc_hd__nand2_1 _18279_ (.A(_02607_),
    .B(_01632_),
    .Y(_02608_));
 sky130_fd_sc_hd__mux2_1 _18280_ (.A0(\core.cpuregs[8][29] ),
    .A1(\core.cpuregs[9][29] ),
    .S(_02404_),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(\core.cpuregs[10][29] ),
    .A1(\core.cpuregs[11][29] ),
    .S(_02406_),
    .X(_02610_));
 sky130_fd_sc_hd__mux2_4 _18282_ (.A0(_02609_),
    .A1(_02610_),
    .S(_10395_),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _18283_ (.A(_02611_),
    .B(_10426_),
    .Y(_02612_));
 sky130_fd_sc_hd__and3_1 _18284_ (.A(_02608_),
    .B(_02612_),
    .C(_02410_),
    .X(_02613_));
 sky130_fd_sc_hd__a31o_1 _18285_ (.A1(_02347_),
    .A2(_02600_),
    .A3(_02604_),
    .B1(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__a21oi_1 _18286_ (.A1(_02614_),
    .A2(_10383_),
    .B1(_10386_),
    .Y(_02615_));
 sky130_fd_sc_hd__mux2_1 _18287_ (.A0(\core.cpuregs[16][29] ),
    .A1(\core.cpuregs[17][29] ),
    .S(_02414_),
    .X(_02616_));
 sky130_fd_sc_hd__mux2_1 _18288_ (.A0(\core.cpuregs[18][29] ),
    .A1(\core.cpuregs[19][29] ),
    .S(_02416_),
    .X(_02617_));
 sky130_fd_sc_hd__mux2_2 _18289_ (.A0(_02616_),
    .A1(_02617_),
    .S(_10344_),
    .X(_02618_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(_02618_),
    .B(_02419_),
    .Y(_02619_));
 sky130_fd_sc_hd__mux2_1 _18291_ (.A0(\core.cpuregs[22][29] ),
    .A1(\core.cpuregs[23][29] ),
    .S(_02421_),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _18292_ (.A0(\core.cpuregs[20][29] ),
    .A1(\core.cpuregs[21][29] ),
    .S(_02423_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _18293_ (.A0(_02620_),
    .A1(_02621_),
    .S(_02425_),
    .X(_02622_));
 sky130_fd_sc_hd__nand2_1 _18294_ (.A(_02622_),
    .B(_10410_),
    .Y(_02623_));
 sky130_fd_sc_hd__mux2_2 _18295_ (.A0(\core.cpuregs[6][29] ),
    .A1(\core.cpuregs[7][29] ),
    .S(_10414_),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(\core.cpuregs[4][29] ),
    .A1(\core.cpuregs[5][29] ),
    .S(_10420_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _18297_ (.A0(_02624_),
    .A1(_02625_),
    .S(_02430_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _18298_ (.A0(\core.cpuregs[0][29] ),
    .A1(\core.cpuregs[1][29] ),
    .S(_10422_),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _18299_ (.A0(\core.cpuregs[2][29] ),
    .A1(\core.cpuregs[3][29] ),
    .S(_10360_),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _18300_ (.A0(_02627_),
    .A1(_02628_),
    .S(_02383_),
    .X(_02629_));
 sky130_fd_sc_hd__and2_1 _18301_ (.A(_02629_),
    .B(_10398_),
    .X(_02630_));
 sky130_fd_sc_hd__a211oi_1 _18302_ (.A1(_10358_),
    .A2(_02626_),
    .B1(_02432_),
    .C1(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__a31o_1 _18303_ (.A1(_02369_),
    .A2(_02619_),
    .A3(_02623_),
    .B1(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_8 _18304_ (.A(_02632_),
    .B(_01746_),
    .Y(_02633_));
 sky130_fd_sc_hd__a22o_1 _18305_ (.A1(\core.decoded_imm[29] ),
    .A2(_04497_),
    .B1(_02615_),
    .B2(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _18306_ (.A0(_02634_),
    .A1(\core.pcpi_rs2[29] ),
    .S(_02441_),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _18307_ (.A(_02635_),
    .X(_00633_));
 sky130_fd_sc_hd__o21ai_2 _18308_ (.A1(_05519_),
    .A2(_04474_),
    .B1(_01649_),
    .Y(_02636_));
 sky130_fd_sc_hd__mux2_1 _18309_ (.A0(\core.cpuregs[16][30] ),
    .A1(\core.cpuregs[17][30] ),
    .S(_01652_),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _18310_ (.A0(\core.cpuregs[18][30] ),
    .A1(\core.cpuregs[19][30] ),
    .S(_01652_),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_1 _18311_ (.A0(_02637_),
    .A1(_02638_),
    .S(_01655_),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_2 _18312_ (.A(_02639_),
    .B(_01657_),
    .Y(_02640_));
 sky130_fd_sc_hd__mux2_1 _18313_ (.A0(\core.cpuregs[22][30] ),
    .A1(\core.cpuregs[23][30] ),
    .S(_01659_),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _18314_ (.A0(\core.cpuregs[20][30] ),
    .A1(\core.cpuregs[21][30] ),
    .S(_01659_),
    .X(_02642_));
 sky130_fd_sc_hd__mux2_1 _18315_ (.A0(_02641_),
    .A1(_02642_),
    .S(_01662_),
    .X(_02643_));
 sky130_fd_sc_hd__nand2_1 _18316_ (.A(_02643_),
    .B(_01664_),
    .Y(_02644_));
 sky130_fd_sc_hd__mux2_1 _18317_ (.A0(\core.cpuregs[6][30] ),
    .A1(\core.cpuregs[7][30] ),
    .S(_01666_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _18318_ (.A0(\core.cpuregs[4][30] ),
    .A1(\core.cpuregs[5][30] ),
    .S(_01666_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _18319_ (.A0(_02645_),
    .A1(_02646_),
    .S(_01662_),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _18320_ (.A0(\core.cpuregs[0][30] ),
    .A1(\core.cpuregs[1][30] ),
    .S(_01671_),
    .X(_02648_));
 sky130_fd_sc_hd__mux2_4 _18321_ (.A0(\core.cpuregs[2][30] ),
    .A1(\core.cpuregs[3][30] ),
    .S(_01671_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _18322_ (.A0(_02648_),
    .A1(_02649_),
    .S(_01674_),
    .X(_02650_));
 sky130_fd_sc_hd__and2_1 _18323_ (.A(_02650_),
    .B(_01676_),
    .X(_02651_));
 sky130_fd_sc_hd__a211oi_2 _18324_ (.A1(_01664_),
    .A2(_02647_),
    .B1(_01651_),
    .C1(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__a31o_1 _18325_ (.A1(_01651_),
    .A2(_02640_),
    .A3(_02644_),
    .B1(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _18326_ (.A0(\core.cpuregs[24][30] ),
    .A1(\core.cpuregs[25][30] ),
    .S(_01681_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _18327_ (.A0(\core.cpuregs[26][30] ),
    .A1(\core.cpuregs[27][30] ),
    .S(_01681_),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _18328_ (.A0(_02654_),
    .A1(_02655_),
    .S(_01655_),
    .X(_02656_));
 sky130_fd_sc_hd__nand2_1 _18329_ (.A(_02656_),
    .B(_01657_),
    .Y(_02657_));
 sky130_fd_sc_hd__mux2_4 _18330_ (.A0(\core.cpuregs[28][30] ),
    .A1(\core.cpuregs[29][30] ),
    .S(_01686_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _18331_ (.A0(\core.cpuregs[30][30] ),
    .A1(\core.cpuregs[31][30] ),
    .S(_01686_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _18332_ (.A0(_02658_),
    .A1(_02659_),
    .S(_01674_),
    .X(_02660_));
 sky130_fd_sc_hd__nand2_1 _18333_ (.A(_02660_),
    .B(_10408_),
    .Y(_02661_));
 sky130_fd_sc_hd__mux2_1 _18334_ (.A0(\core.cpuregs[8][30] ),
    .A1(\core.cpuregs[9][30] ),
    .S(_01691_),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _18335_ (.A0(\core.cpuregs[10][30] ),
    .A1(\core.cpuregs[11][30] ),
    .S(_01691_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _18336_ (.A0(_02662_),
    .A1(_02663_),
    .S(_10396_),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _18337_ (.A0(\core.cpuregs[12][30] ),
    .A1(\core.cpuregs[13][30] ),
    .S(_01695_),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _18338_ (.A0(\core.cpuregs[14][30] ),
    .A1(\core.cpuregs[15][30] ),
    .S(_10350_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _18339_ (.A0(_02665_),
    .A1(_02666_),
    .S(_01698_),
    .X(_02667_));
 sky130_fd_sc_hd__and2_1 _18340_ (.A(_02667_),
    .B(_10369_),
    .X(_02668_));
 sky130_fd_sc_hd__a211oi_1 _18341_ (.A1(_01676_),
    .A2(_02664_),
    .B1(_01680_),
    .C1(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a31o_1 _18342_ (.A1(_01680_),
    .A2(_02657_),
    .A3(_02661_),
    .B1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__a21oi_2 _18343_ (.A1(_02670_),
    .A2(_10384_),
    .B1(_10387_),
    .Y(_02671_));
 sky130_fd_sc_hd__a21boi_1 _18344_ (.A1(_10431_),
    .A2(_02653_),
    .B1_N(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__o22a_1 _18345_ (.A1(\core.pcpi_rs2[30] ),
    .A2(_01649_),
    .B1(_02636_),
    .B2(_02672_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _18346_ (.A0(\core.cpuregs[24][31] ),
    .A1(\core.cpuregs[25][31] ),
    .S(_10342_),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _18347_ (.A0(\core.cpuregs[26][31] ),
    .A1(\core.cpuregs[27][31] ),
    .S(_01695_),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _18348_ (.A0(_02673_),
    .A1(_02674_),
    .S(_01698_),
    .X(_02675_));
 sky130_fd_sc_hd__nand2_1 _18349_ (.A(_02675_),
    .B(_10399_),
    .Y(_02676_));
 sky130_fd_sc_hd__mux2_1 _18350_ (.A0(\core.cpuregs[28][31] ),
    .A1(\core.cpuregs[29][31] ),
    .S(_10353_),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _18351_ (.A0(\core.cpuregs[30][31] ),
    .A1(\core.cpuregs[31][31] ),
    .S(_10411_),
    .X(_02678_));
 sky130_fd_sc_hd__mux2_1 _18352_ (.A0(_02677_),
    .A1(_02678_),
    .S(_02397_),
    .X(_02679_));
 sky130_fd_sc_hd__nand2_1 _18353_ (.A(_02679_),
    .B(_01700_),
    .Y(_02680_));
 sky130_fd_sc_hd__mux2_1 _18354_ (.A0(\core.cpuregs[12][31] ),
    .A1(\core.cpuregs[13][31] ),
    .S(_10363_),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _18355_ (.A0(\core.cpuregs[14][31] ),
    .A1(\core.cpuregs[15][31] ),
    .S(_01670_),
    .X(_02682_));
 sky130_fd_sc_hd__mux2_1 _18356_ (.A0(_02681_),
    .A1(_02682_),
    .S(_10376_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _18357_ (.A(_02683_),
    .B(_01632_),
    .Y(_02684_));
 sky130_fd_sc_hd__mux2_1 _18358_ (.A0(\core.cpuregs[8][31] ),
    .A1(\core.cpuregs[9][31] ),
    .S(_02404_),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _18359_ (.A0(\core.cpuregs[10][31] ),
    .A1(\core.cpuregs[11][31] ),
    .S(_02406_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _18360_ (.A0(_02685_),
    .A1(_02686_),
    .S(_10395_),
    .X(_02687_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(_02687_),
    .B(_10426_),
    .Y(_02688_));
 sky130_fd_sc_hd__and3_1 _18362_ (.A(_02684_),
    .B(_02688_),
    .C(_02410_),
    .X(_02689_));
 sky130_fd_sc_hd__a31o_1 _18363_ (.A1(_04573_),
    .A2(_02676_),
    .A3(_02680_),
    .B1(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__a21oi_2 _18364_ (.A1(_02690_),
    .A2(_10383_),
    .B1(_10386_),
    .Y(_02691_));
 sky130_fd_sc_hd__mux2_1 _18365_ (.A0(\core.cpuregs[16][31] ),
    .A1(\core.cpuregs[17][31] ),
    .S(_02414_),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _18366_ (.A0(\core.cpuregs[18][31] ),
    .A1(\core.cpuregs[19][31] ),
    .S(_02416_),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_4 _18367_ (.A0(_02692_),
    .A1(_02693_),
    .S(_10344_),
    .X(_02694_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(_02694_),
    .B(_02419_),
    .Y(_02695_));
 sky130_fd_sc_hd__mux2_1 _18369_ (.A0(\core.cpuregs[22][31] ),
    .A1(\core.cpuregs[23][31] ),
    .S(_02421_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _18370_ (.A0(\core.cpuregs[20][31] ),
    .A1(\core.cpuregs[21][31] ),
    .S(_02423_),
    .X(_02697_));
 sky130_fd_sc_hd__mux2_4 _18371_ (.A0(_02696_),
    .A1(_02697_),
    .S(_02425_),
    .X(_02698_));
 sky130_fd_sc_hd__nand2_1 _18372_ (.A(_02698_),
    .B(_10410_),
    .Y(_02699_));
 sky130_fd_sc_hd__mux2_1 _18373_ (.A0(\core.cpuregs[6][31] ),
    .A1(\core.cpuregs[7][31] ),
    .S(_10414_),
    .X(_02700_));
 sky130_fd_sc_hd__mux2_1 _18374_ (.A0(\core.cpuregs[4][31] ),
    .A1(\core.cpuregs[5][31] ),
    .S(_10420_),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _18375_ (.A0(_02700_),
    .A1(_02701_),
    .S(_02430_),
    .X(_02702_));
 sky130_fd_sc_hd__mux2_1 _18376_ (.A0(\core.cpuregs[0][31] ),
    .A1(\core.cpuregs[1][31] ),
    .S(_10422_),
    .X(_02703_));
 sky130_fd_sc_hd__mux2_1 _18377_ (.A0(\core.cpuregs[2][31] ),
    .A1(\core.cpuregs[3][31] ),
    .S(_10360_),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _18378_ (.A0(_02703_),
    .A1(_02704_),
    .S(_10366_),
    .X(_02705_));
 sky130_fd_sc_hd__and2_1 _18379_ (.A(_02705_),
    .B(_10398_),
    .X(_02706_));
 sky130_fd_sc_hd__a211oi_1 _18380_ (.A1(_10358_),
    .A2(_02702_),
    .B1(_02432_),
    .C1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a31o_1 _18381_ (.A1(_10337_),
    .A2(_02695_),
    .A3(_02699_),
    .B1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(_02708_),
    .B(_01746_),
    .Y(_02709_));
 sky130_fd_sc_hd__a22o_1 _18383_ (.A1(\core.decoded_imm[31] ),
    .A2(_04497_),
    .B1(_02691_),
    .B2(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _18384_ (.A0(_02710_),
    .A1(\core.pcpi_rs2[31] ),
    .S(_02441_),
    .X(_02711_));
 sky130_fd_sc_hd__buf_1 _18385_ (.A(_02711_),
    .X(_00635_));
 sky130_fd_sc_hd__o22a_1 _18386_ (.A1(_04435_),
    .A2(_10055_),
    .B1(_10056_),
    .B2(_10248_),
    .X(_02712_));
 sky130_fd_sc_hd__nor2_4 _18387_ (.A(_06372_),
    .B(_02712_),
    .Y(_00636_));
 sky130_fd_sc_hd__o2bb2a_1 _18388_ (.A1_N(\core.instr_bltu ),
    .A2_N(_10226_),
    .B1(_10056_),
    .B2(_10229_),
    .X(_02713_));
 sky130_fd_sc_hd__nor2_1 _18389_ (.A(_06372_),
    .B(_02713_),
    .Y(_00637_));
 sky130_fd_sc_hd__mux2_1 _18390_ (.A0(net5),
    .A1(\core.mem_rdata_q[13] ),
    .S(_05923_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _18391_ (.A(_02714_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _18392_ (.A0(net6),
    .A1(\core.mem_rdata_q[14] ),
    .S(_05923_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_2 _18393_ (.A(_02715_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _18394_ (.A0(net4),
    .A1(\core.mem_rdata_q[12] ),
    .S(_05940_),
    .X(_02716_));
 sky130_fd_sc_hd__clkbuf_1 _18395_ (.A(_02716_),
    .X(_01355_));
 sky130_fd_sc_hd__nor3_1 _18396_ (.A(_01356_),
    .B(_01357_),
    .C(_01355_),
    .Y(_02717_));
 sky130_fd_sc_hd__and3_1 _18397_ (.A(_10031_),
    .B(_10150_),
    .C(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_4 _18398_ (.A(_05932_),
    .X(_02719_));
 sky130_fd_sc_hd__mux2_1 _18399_ (.A0(_02718_),
    .A1(\core.instr_jalr ),
    .S(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_1 _18400_ (.A(_02720_),
    .X(_00638_));
 sky130_fd_sc_hd__nand2_2 _18401_ (.A(_10055_),
    .B(\core.is_lb_lh_lw_lbu_lhu ),
    .Y(_02721_));
 sky130_fd_sc_hd__inv_2 _18402_ (.A(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__a22o_1 _18403_ (.A1(\core.instr_lb ),
    .A2(_10218_),
    .B1(_10155_),
    .B2(_02722_),
    .X(_00639_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(_09327_),
    .B(_09950_),
    .Y(_02723_));
 sky130_fd_sc_hd__clkbuf_4 _18405_ (.A(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_2 _18406_ (.A(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_8 _18407_ (.A0(\core.cpuregs[20][0] ),
    .A1(_10062_),
    .S(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_1 _18408_ (.A(_02726_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(\core.cpuregs[20][1] ),
    .A1(_10069_),
    .S(_02725_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _18410_ (.A(_02727_),
    .X(_00641_));
 sky130_fd_sc_hd__buf_2 _18411_ (.A(_02724_),
    .X(_02728_));
 sky130_fd_sc_hd__mux2_2 _18412_ (.A0(\core.cpuregs[20][2] ),
    .A1(_10071_),
    .S(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__buf_1 _18413_ (.A(_02729_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _18414_ (.A0(\core.cpuregs[20][3] ),
    .A1(_10074_),
    .S(_02728_),
    .X(_02730_));
 sky130_fd_sc_hd__buf_1 _18415_ (.A(_02730_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(\core.cpuregs[20][4] ),
    .A1(_10076_),
    .S(_02728_),
    .X(_02731_));
 sky130_fd_sc_hd__buf_1 _18417_ (.A(_02731_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _18418_ (.A0(\core.cpuregs[20][5] ),
    .A1(_10078_),
    .S(_02728_),
    .X(_02732_));
 sky130_fd_sc_hd__buf_1 _18419_ (.A(_02732_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _18420_ (.A0(\core.cpuregs[20][6] ),
    .A1(_10080_),
    .S(_02728_),
    .X(_02733_));
 sky130_fd_sc_hd__clkbuf_1 _18421_ (.A(_02733_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _18422_ (.A0(\core.cpuregs[20][7] ),
    .A1(_10082_),
    .S(_02728_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _18423_ (.A(_02734_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18424_ (.A0(\core.cpuregs[20][8] ),
    .A1(_10084_),
    .S(_02724_),
    .X(_02735_));
 sky130_fd_sc_hd__clkbuf_1 _18425_ (.A(_02735_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_2 _18426_ (.A0(\core.cpuregs[20][9] ),
    .A1(_10086_),
    .S(_02724_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_1 _18427_ (.A(_02736_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18428_ (.A0(\core.cpuregs[20][10] ),
    .A1(_10088_),
    .S(_02724_),
    .X(_02737_));
 sky130_fd_sc_hd__clkbuf_1 _18429_ (.A(_02737_),
    .X(_00650_));
 sky130_fd_sc_hd__inv_2 _18430_ (.A(_02723_),
    .Y(_02738_));
 sky130_fd_sc_hd__clkbuf_2 _18431_ (.A(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _18432_ (.A0(_10090_),
    .A1(\core.cpuregs[20][11] ),
    .S(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__clkbuf_1 _18433_ (.A(_02740_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18434_ (.A0(\core.cpuregs[20][12] ),
    .A1(_10094_),
    .S(_02724_),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_1 _18435_ (.A(_02741_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_2 _18436_ (.A0(_10096_),
    .A1(\core.cpuregs[20][13] ),
    .S(_02739_),
    .X(_02742_));
 sky130_fd_sc_hd__buf_1 _18437_ (.A(_02742_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18438_ (.A0(_10098_),
    .A1(\core.cpuregs[20][14] ),
    .S(_02738_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _18439_ (.A(_02743_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18440_ (.A0(_10100_),
    .A1(\core.cpuregs[20][15] ),
    .S(_02738_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_1 _18441_ (.A(_02744_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_4 _18442_ (.A0(_10102_),
    .A1(\core.cpuregs[20][16] ),
    .S(_02738_),
    .X(_02745_));
 sky130_fd_sc_hd__buf_1 _18443_ (.A(_02745_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18444_ (.A0(_10104_),
    .A1(\core.cpuregs[20][17] ),
    .S(_02738_),
    .X(_02746_));
 sky130_fd_sc_hd__clkbuf_1 _18445_ (.A(_02746_),
    .X(_00657_));
 sky130_fd_sc_hd__nand2_1 _18446_ (.A(_02739_),
    .B(\core.cpuregs[20][18] ),
    .Y(_02747_));
 sky130_fd_sc_hd__a21bo_1 _18447_ (.A1(_09837_),
    .A2(_02725_),
    .B1_N(_02747_),
    .X(_00658_));
 sky130_fd_sc_hd__clkbuf_4 _18448_ (.A(_02725_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_1 _18449_ (.A(_10107_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__clkbuf_4 _18450_ (.A(_02739_),
    .X(_02750_));
 sky130_fd_sc_hd__nand2_2 _18451_ (.A(_02750_),
    .B(\core.cpuregs[20][19] ),
    .Y(_02751_));
 sky130_fd_sc_hd__nand2_1 _18452_ (.A(_02749_),
    .B(_02751_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_10112_),
    .B(_02748_),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_2 _18454_ (.A(_02750_),
    .B(\core.cpuregs[20][20] ),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _18455_ (.A(_02752_),
    .B(_02753_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_1 _18456_ (.A(_10115_),
    .B(_02748_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _18457_ (.A(_02750_),
    .B(\core.cpuregs[20][21] ),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _18458_ (.A(_02754_),
    .B(_02755_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _18459_ (.A(_10118_),
    .B(_02748_),
    .Y(_02756_));
 sky130_fd_sc_hd__nand2_1 _18460_ (.A(_02750_),
    .B(\core.cpuregs[20][22] ),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _18461_ (.A(_02756_),
    .B(_02757_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _18462_ (.A(_10121_),
    .B(_02748_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_02750_),
    .B(\core.cpuregs[20][23] ),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2_1 _18464_ (.A(_02758_),
    .B(_02759_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _18465_ (.A(_10124_),
    .B(_02748_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _18466_ (.A(_02750_),
    .B(\core.cpuregs[20][24] ),
    .Y(_02761_));
 sky130_fd_sc_hd__nand2_1 _18467_ (.A(_02760_),
    .B(_02761_),
    .Y(_00664_));
 sky130_fd_sc_hd__clkbuf_2 _18468_ (.A(_02725_),
    .X(_02762_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(_10127_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__buf_2 _18470_ (.A(_02739_),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_4 _18471_ (.A(_02764_),
    .B(\core.cpuregs[20][25] ),
    .Y(_02765_));
 sky130_fd_sc_hd__nand2_1 _18472_ (.A(_02763_),
    .B(_02765_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _18473_ (.A(_10132_),
    .B(_02762_),
    .Y(_02766_));
 sky130_fd_sc_hd__nand2_1 _18474_ (.A(_02764_),
    .B(net195),
    .Y(_02767_));
 sky130_fd_sc_hd__nand2_1 _18475_ (.A(_02766_),
    .B(_02767_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_2 _18476_ (.A(_10135_),
    .B(_02762_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_4 _18477_ (.A(_02764_),
    .B(\core.cpuregs[20][27] ),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_1 _18478_ (.A(_02768_),
    .B(_02769_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_2 _18479_ (.A(_10138_),
    .B(_02762_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_2 _18480_ (.A(_02764_),
    .B(\core.cpuregs[20][28] ),
    .Y(_02771_));
 sky130_fd_sc_hd__nand2_1 _18481_ (.A(_02770_),
    .B(_02771_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(_10141_),
    .B(_02762_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _18483_ (.A(_02764_),
    .B(\core.cpuregs[20][29] ),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_1 _18484_ (.A(_02772_),
    .B(_02773_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_2 _18485_ (.A(_10144_),
    .B(_02762_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _18486_ (.A(_02764_),
    .B(\core.cpuregs[20][30] ),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_02774_),
    .B(_02775_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_10147_),
    .B(_02725_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_02739_),
    .B(\core.cpuregs[20][31] ),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _18490_ (.A(_02776_),
    .B(_02777_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _18491_ (.A(_09324_),
    .B(_10064_),
    .Y(_02778_));
 sky130_fd_sc_hd__nor2_1 _18492_ (.A(_09811_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__clkbuf_2 _18493_ (.A(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_2 _18494_ (.A(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_2 _18495_ (.A0(\core.cpuregs[25][0] ),
    .A1(_10062_),
    .S(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_2 _18496_ (.A(_02782_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_4 _18497_ (.A0(\core.cpuregs[25][1] ),
    .A1(_10069_),
    .S(_02781_),
    .X(_02783_));
 sky130_fd_sc_hd__clkbuf_1 _18498_ (.A(_02783_),
    .X(_00673_));
 sky130_fd_sc_hd__clkbuf_4 _18499_ (.A(_02780_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _18500_ (.A0(\core.cpuregs[25][2] ),
    .A1(_10071_),
    .S(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_1 _18501_ (.A(_02785_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18502_ (.A0(\core.cpuregs[25][3] ),
    .A1(_10074_),
    .S(_02784_),
    .X(_02786_));
 sky130_fd_sc_hd__buf_1 _18503_ (.A(_02786_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _18504_ (.A0(\core.cpuregs[25][4] ),
    .A1(_10076_),
    .S(_02784_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _18505_ (.A(_02787_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18506_ (.A0(\core.cpuregs[25][5] ),
    .A1(_10078_),
    .S(_02784_),
    .X(_02788_));
 sky130_fd_sc_hd__buf_1 _18507_ (.A(_02788_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _18508_ (.A0(\core.cpuregs[25][6] ),
    .A1(_10080_),
    .S(_02784_),
    .X(_02789_));
 sky130_fd_sc_hd__buf_1 _18509_ (.A(_02789_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _18510_ (.A0(\core.cpuregs[25][7] ),
    .A1(_10082_),
    .S(_02784_),
    .X(_02790_));
 sky130_fd_sc_hd__clkbuf_1 _18511_ (.A(_02790_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _18512_ (.A0(\core.cpuregs[25][8] ),
    .A1(_10084_),
    .S(_02780_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _18513_ (.A(_02791_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _18514_ (.A0(\core.cpuregs[25][9] ),
    .A1(_10086_),
    .S(_02780_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _18515_ (.A(_02792_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18516_ (.A0(\core.cpuregs[25][10] ),
    .A1(_10088_),
    .S(_02780_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_1 _18517_ (.A(_02793_),
    .X(_00682_));
 sky130_fd_sc_hd__inv_2 _18518_ (.A(_02779_),
    .Y(_02794_));
 sky130_fd_sc_hd__clkbuf_2 _18519_ (.A(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _18520_ (.A0(_10090_),
    .A1(\core.cpuregs[25][11] ),
    .S(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__buf_1 _18521_ (.A(_02796_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _18522_ (.A0(\core.cpuregs[25][12] ),
    .A1(_10094_),
    .S(_02780_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_1 _18523_ (.A(_02797_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _18524_ (.A0(_10096_),
    .A1(\core.cpuregs[25][13] ),
    .S(_02795_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _18525_ (.A(_02798_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _18526_ (.A0(_10098_),
    .A1(\core.cpuregs[25][14] ),
    .S(_02794_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _18527_ (.A(_02799_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _18528_ (.A0(_10100_),
    .A1(\core.cpuregs[25][15] ),
    .S(_02794_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_1 _18529_ (.A(_02800_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _18530_ (.A0(_10102_),
    .A1(\core.cpuregs[25][16] ),
    .S(_02794_),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_1 _18531_ (.A(_02801_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _18532_ (.A0(_10104_),
    .A1(\core.cpuregs[25][17] ),
    .S(_02794_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _18533_ (.A(_02802_),
    .X(_00689_));
 sky130_fd_sc_hd__nand2_1 _18534_ (.A(_02795_),
    .B(\core.cpuregs[25][18] ),
    .Y(_02803_));
 sky130_fd_sc_hd__a21bo_1 _18535_ (.A1(_09837_),
    .A2(_02781_),
    .B1_N(_02803_),
    .X(_00690_));
 sky130_fd_sc_hd__clkbuf_2 _18536_ (.A(_02781_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_1 _18537_ (.A(_10107_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18538_ (.A(_02795_),
    .X(_02806_));
 sky130_fd_sc_hd__nand2_1 _18539_ (.A(_02806_),
    .B(\core.cpuregs[25][19] ),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _18540_ (.A(_02805_),
    .B(_02807_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_2 _18541_ (.A(_10112_),
    .B(_02804_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _18542_ (.A(_02806_),
    .B(\core.cpuregs[25][20] ),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(_02808_),
    .B(_02809_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _18544_ (.A(_10115_),
    .B(_02804_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2_1 _18545_ (.A(_02806_),
    .B(\core.cpuregs[25][21] ),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _18546_ (.A(_02810_),
    .B(_02811_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(_10118_),
    .B(_02804_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _18548_ (.A(_02806_),
    .B(\core.cpuregs[25][22] ),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_1 _18549_ (.A(_02812_),
    .B(_02813_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_2 _18550_ (.A(_10121_),
    .B(_02804_),
    .Y(_02814_));
 sky130_fd_sc_hd__nand2_1 _18551_ (.A(_02806_),
    .B(\core.cpuregs[25][23] ),
    .Y(_02815_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(_02814_),
    .B(_02815_),
    .Y(_00695_));
 sky130_fd_sc_hd__nand2_1 _18553_ (.A(_10124_),
    .B(_02804_),
    .Y(_02816_));
 sky130_fd_sc_hd__nand2_1 _18554_ (.A(_02806_),
    .B(\core.cpuregs[25][24] ),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _18555_ (.A(_02816_),
    .B(_02817_),
    .Y(_00696_));
 sky130_fd_sc_hd__clkbuf_4 _18556_ (.A(_02781_),
    .X(_02818_));
 sky130_fd_sc_hd__nand2_1 _18557_ (.A(_10127_),
    .B(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18558_ (.A(_02795_),
    .X(_02820_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(_02820_),
    .B(\core.cpuregs[25][25] ),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(_02819_),
    .B(_02821_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _18561_ (.A(_10132_),
    .B(_02818_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _18562_ (.A(_02820_),
    .B(\core.cpuregs[25][26] ),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _18563_ (.A(_02822_),
    .B(_02823_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _18564_ (.A(_10135_),
    .B(_02818_),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _18565_ (.A(_02820_),
    .B(\core.cpuregs[25][27] ),
    .Y(_02825_));
 sky130_fd_sc_hd__nand2_1 _18566_ (.A(_02824_),
    .B(_02825_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(_10138_),
    .B(_02818_),
    .Y(_02826_));
 sky130_fd_sc_hd__nand2_1 _18568_ (.A(_02820_),
    .B(\core.cpuregs[25][28] ),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(_02826_),
    .B(_02827_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _18570_ (.A(_10141_),
    .B(_02818_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(_02820_),
    .B(\core.cpuregs[25][29] ),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _18572_ (.A(_02828_),
    .B(_02829_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_2 _18573_ (.A(_10144_),
    .B(_02818_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(_02820_),
    .B(\core.cpuregs[25][30] ),
    .Y(_02831_));
 sky130_fd_sc_hd__nand2_1 _18575_ (.A(_02830_),
    .B(_02831_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _18576_ (.A(_10147_),
    .B(_02781_),
    .Y(_02832_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(_02795_),
    .B(\core.cpuregs[25][31] ),
    .Y(_02833_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(_02832_),
    .B(_02833_),
    .Y(_00703_));
 sky130_fd_sc_hd__and3_1 _18579_ (.A(_09554_),
    .B(_09320_),
    .C(_10064_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_2 _18580_ (.A(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_4 _18581_ (.A(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _18582_ (.A0(\core.cpuregs[1][0] ),
    .A1(_10062_),
    .S(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_8 _18583_ (.A(_02837_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18584_ (.A0(\core.cpuregs[1][1] ),
    .A1(_10069_),
    .S(_02836_),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _18585_ (.A(_02838_),
    .X(_00705_));
 sky130_fd_sc_hd__clkbuf_4 _18586_ (.A(_02835_),
    .X(_02839_));
 sky130_fd_sc_hd__mux2_1 _18587_ (.A0(\core.cpuregs[1][2] ),
    .A1(_10071_),
    .S(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _18588_ (.A(_02840_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _18589_ (.A0(\core.cpuregs[1][3] ),
    .A1(_10074_),
    .S(_02839_),
    .X(_02841_));
 sky130_fd_sc_hd__buf_1 _18590_ (.A(_02841_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _18591_ (.A0(\core.cpuregs[1][4] ),
    .A1(_10076_),
    .S(_02839_),
    .X(_02842_));
 sky130_fd_sc_hd__buf_1 _18592_ (.A(_02842_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _18593_ (.A0(\core.cpuregs[1][5] ),
    .A1(_10078_),
    .S(_02839_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _18594_ (.A(_02843_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _18595_ (.A0(\core.cpuregs[1][6] ),
    .A1(_10080_),
    .S(_02839_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _18596_ (.A(_02844_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _18597_ (.A0(\core.cpuregs[1][7] ),
    .A1(_10082_),
    .S(_02839_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _18598_ (.A(_02845_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _18599_ (.A0(\core.cpuregs[1][8] ),
    .A1(_10084_),
    .S(_02835_),
    .X(_02846_));
 sky130_fd_sc_hd__buf_1 _18600_ (.A(_02846_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _18601_ (.A0(\core.cpuregs[1][9] ),
    .A1(_10086_),
    .S(_02835_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _18602_ (.A(_02847_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _18603_ (.A0(\core.cpuregs[1][10] ),
    .A1(_10088_),
    .S(_02835_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _18604_ (.A(_02848_),
    .X(_00714_));
 sky130_fd_sc_hd__inv_2 _18605_ (.A(_02834_),
    .Y(_02849_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18606_ (.A(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _18607_ (.A0(_10090_),
    .A1(\core.cpuregs[1][11] ),
    .S(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _18608_ (.A(_02851_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _18609_ (.A0(\core.cpuregs[1][12] ),
    .A1(_10094_),
    .S(_02835_),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _18610_ (.A(_02852_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _18611_ (.A0(_10096_),
    .A1(\core.cpuregs[1][13] ),
    .S(_02850_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _18612_ (.A(_02853_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _18613_ (.A0(_10098_),
    .A1(\core.cpuregs[1][14] ),
    .S(_02849_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _18614_ (.A(_02854_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_2 _18615_ (.A0(_10100_),
    .A1(\core.cpuregs[1][15] ),
    .S(_02849_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _18616_ (.A(_02855_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _18617_ (.A0(_10102_),
    .A1(\core.cpuregs[1][16] ),
    .S(_02849_),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _18618_ (.A(_02856_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _18619_ (.A0(_10104_),
    .A1(\core.cpuregs[1][17] ),
    .S(_02849_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _18620_ (.A(_02857_),
    .X(_00721_));
 sky130_fd_sc_hd__and2_1 _18621_ (.A(_02850_),
    .B(\core.cpuregs[1][18] ),
    .X(_02858_));
 sky130_fd_sc_hd__a21o_1 _18622_ (.A1(_09779_),
    .A2(_02836_),
    .B1(_02858_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_2 _18623_ (.A(_02836_),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(_10107_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__buf_4 _18625_ (.A(_02850_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_1 _18626_ (.A(_02861_),
    .B(\core.cpuregs[1][19] ),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _18627_ (.A(_02860_),
    .B(_02862_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _18628_ (.A(_10112_),
    .B(_02859_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_1 _18629_ (.A(_02861_),
    .B(\core.cpuregs[1][20] ),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _18630_ (.A(_02863_),
    .B(_02864_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _18631_ (.A(_10115_),
    .B(_02859_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(_02861_),
    .B(net145),
    .Y(_02866_));
 sky130_fd_sc_hd__nand2_1 _18633_ (.A(_02865_),
    .B(_02866_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_1 _18634_ (.A(_10118_),
    .B(_02859_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_1 _18635_ (.A(_02861_),
    .B(\core.cpuregs[1][22] ),
    .Y(_02868_));
 sky130_fd_sc_hd__nand2_1 _18636_ (.A(_02867_),
    .B(_02868_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_1 _18637_ (.A(_10121_),
    .B(_02859_),
    .Y(_02869_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(_02861_),
    .B(\core.cpuregs[1][23] ),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(_02869_),
    .B(_02870_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_1 _18640_ (.A(_10124_),
    .B(_02859_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(_02861_),
    .B(\core.cpuregs[1][24] ),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(_02871_),
    .B(_02872_),
    .Y(_00728_));
 sky130_fd_sc_hd__buf_4 _18643_ (.A(_02836_),
    .X(_02873_));
 sky130_fd_sc_hd__nand2_4 _18644_ (.A(_10127_),
    .B(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__clkbuf_2 _18645_ (.A(_02850_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_2 _18646_ (.A(_02875_),
    .B(\core.cpuregs[1][25] ),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(_02874_),
    .B(_02876_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _18648_ (.A(_10132_),
    .B(_02873_),
    .Y(_02877_));
 sky130_fd_sc_hd__nand2_1 _18649_ (.A(_02875_),
    .B(\core.cpuregs[1][26] ),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _18650_ (.A(_02877_),
    .B(_02878_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _18651_ (.A(_10135_),
    .B(_02873_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_4 _18652_ (.A(_02875_),
    .B(\core.cpuregs[1][27] ),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _18653_ (.A(_02879_),
    .B(_02880_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(_10138_),
    .B(_02873_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _18655_ (.A(_02875_),
    .B(\core.cpuregs[1][28] ),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_1 _18656_ (.A(_02881_),
    .B(_02882_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_2 _18657_ (.A(_10141_),
    .B(_02873_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_2 _18658_ (.A(_02875_),
    .B(\core.cpuregs[1][29] ),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _18659_ (.A(_02883_),
    .B(_02884_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _18660_ (.A(_10144_),
    .B(_02873_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _18661_ (.A(_02875_),
    .B(net128),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_1 _18662_ (.A(_02885_),
    .B(_02886_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _18663_ (.A(_10147_),
    .B(_02836_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand2_1 _18664_ (.A(_02850_),
    .B(\core.cpuregs[1][31] ),
    .Y(_02888_));
 sky130_fd_sc_hd__nand2_1 _18665_ (.A(_02887_),
    .B(_02888_),
    .Y(_00735_));
 sky130_fd_sc_hd__clkbuf_2 _18666_ (.A(_05940_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _18667_ (.A0(net30),
    .A1(\core.mem_rdata_q[7] ),
    .S(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_1 _18668_ (.A(_02890_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _18669_ (.A0(_01350_),
    .A1(\core.decoded_rd[0] ),
    .S(_02719_),
    .X(_02891_));
 sky130_fd_sc_hd__buf_1 _18670_ (.A(_02891_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _18671_ (.A0(net31),
    .A1(\core.mem_rdata_q[8] ),
    .S(_02889_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_2 _18672_ (.A(_02892_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _18673_ (.A0(_01351_),
    .A1(\core.decoded_rd[1] ),
    .S(_02719_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_1 _18674_ (.A(_02893_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _18675_ (.A0(net32),
    .A1(\core.mem_rdata_q[9] ),
    .S(_02889_),
    .X(_02894_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18676_ (.A(_02894_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _18677_ (.A0(_01352_),
    .A1(\core.decoded_rd[2] ),
    .S(_02719_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _18678_ (.A(_02895_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _18679_ (.A0(net2),
    .A1(\core.mem_rdata_q[10] ),
    .S(_02889_),
    .X(_02896_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18680_ (.A(_02896_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _18681_ (.A0(_01353_),
    .A1(\core.decoded_rd[3] ),
    .S(_02719_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _18682_ (.A(_02897_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _18683_ (.A0(net3),
    .A1(\core.mem_rdata_q[11] ),
    .S(_02889_),
    .X(_02898_));
 sky130_fd_sc_hd__buf_1 _18684_ (.A(_02898_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _18685_ (.A0(_01354_),
    .A1(\core.decoded_rd[4] ),
    .S(_02719_),
    .X(_02899_));
 sky130_fd_sc_hd__buf_1 _18686_ (.A(_02899_),
    .X(_00740_));
 sky130_fd_sc_hd__or3_1 _18687_ (.A(\core.instr_jalr ),
    .B(\core.is_lb_lh_lw_lbu_lhu ),
    .C(\core.is_alu_reg_imm ),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_4 _18688_ (.A(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__a22o_1 _18689_ (.A1(_04468_),
    .A2(\core.mem_rdata_q[7] ),
    .B1(_02901_),
    .B2(\core.mem_rdata_q[20] ),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_4 _18690_ (.A(_10215_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _18691_ (.A0(_02902_),
    .A1(\core.decoded_imm[0] ),
    .S(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__buf_1 _18692_ (.A(_02904_),
    .X(_00741_));
 sky130_fd_sc_hd__buf_4 _18693_ (.A(_05932_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _18694_ (.A0(_01364_),
    .A1(_05942_),
    .S(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__buf_1 _18695_ (.A(_02906_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _18696_ (.A0(_01365_),
    .A1(\core.decoded_imm_j[2] ),
    .S(_02905_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_1 _18697_ (.A(_02907_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_8 _18698_ (.A0(_01366_),
    .A1(_04575_),
    .S(_02905_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _18699_ (.A(_02908_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _18700_ (.A0(_01367_),
    .A1(_04576_),
    .S(_02905_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _18701_ (.A(_02909_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _18702_ (.A0(net18),
    .A1(\core.mem_rdata_q[25] ),
    .S(_02889_),
    .X(_02910_));
 sky130_fd_sc_hd__buf_1 _18703_ (.A(_02910_),
    .X(_01368_));
 sky130_fd_sc_hd__buf_4 _18704_ (.A(_05932_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _18705_ (.A0(_01368_),
    .A1(\core.decoded_imm_j[5] ),
    .S(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_1 _18706_ (.A(_02912_),
    .X(_00746_));
 sky130_fd_sc_hd__buf_4 _18707_ (.A(_05923_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _18708_ (.A0(net19),
    .A1(\core.mem_rdata_q[26] ),
    .S(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_2 _18709_ (.A(_02914_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _18710_ (.A0(_01369_),
    .A1(\core.decoded_imm_j[6] ),
    .S(_02911_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _18711_ (.A(_02915_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _18712_ (.A0(net20),
    .A1(\core.mem_rdata_q[27] ),
    .S(_02913_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _18713_ (.A(_02916_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _18714_ (.A0(_01370_),
    .A1(\core.decoded_imm_j[7] ),
    .S(_02911_),
    .X(_02917_));
 sky130_fd_sc_hd__buf_1 _18715_ (.A(_02917_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _18716_ (.A0(net21),
    .A1(\core.mem_rdata_q[28] ),
    .S(_02913_),
    .X(_02918_));
 sky130_fd_sc_hd__buf_1 _18717_ (.A(_02918_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _18718_ (.A0(_01371_),
    .A1(\core.decoded_imm_j[8] ),
    .S(_02911_),
    .X(_02919_));
 sky130_fd_sc_hd__buf_1 _18719_ (.A(_02919_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _18720_ (.A0(net22),
    .A1(\core.mem_rdata_q[29] ),
    .S(_02913_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _18721_ (.A(_02920_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _18722_ (.A0(_01372_),
    .A1(\core.decoded_imm_j[9] ),
    .S(_02911_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_4 _18723_ (.A(_02921_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _18724_ (.A0(net24),
    .A1(\core.mem_rdata_q[30] ),
    .S(_02913_),
    .X(_02922_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18725_ (.A(_02922_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _18726_ (.A0(_01373_),
    .A1(\core.decoded_imm_j[10] ),
    .S(_02911_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_4 _18727_ (.A(_02923_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _18728_ (.A0(_01363_),
    .A1(_04577_),
    .S(_02905_),
    .X(_02924_));
 sky130_fd_sc_hd__buf_1 _18729_ (.A(_02924_),
    .X(_00752_));
 sky130_fd_sc_hd__clkbuf_2 _18730_ (.A(_05932_),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _18731_ (.A0(_01355_),
    .A1(\core.decoded_imm_j[12] ),
    .S(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__buf_1 _18732_ (.A(_02926_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _18733_ (.A0(_01356_),
    .A1(\core.decoded_imm_j[13] ),
    .S(_02925_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _18734_ (.A(_02927_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _18735_ (.A0(_01357_),
    .A1(\core.decoded_imm_j[14] ),
    .S(_02925_),
    .X(_02928_));
 sky130_fd_sc_hd__buf_1 _18736_ (.A(_02928_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _18737_ (.A0(_01358_),
    .A1(\core.decoded_imm_j[15] ),
    .S(_02905_),
    .X(_02929_));
 sky130_fd_sc_hd__buf_1 _18738_ (.A(_02929_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _18739_ (.A0(_01359_),
    .A1(\core.decoded_imm_j[16] ),
    .S(_04978_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _18740_ (.A(_02930_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _18741_ (.A0(_01360_),
    .A1(\core.decoded_imm_j[17] ),
    .S(_04978_),
    .X(_02931_));
 sky130_fd_sc_hd__buf_1 _18742_ (.A(_02931_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _18743_ (.A0(_01361_),
    .A1(\core.decoded_imm_j[18] ),
    .S(_04978_),
    .X(_02932_));
 sky130_fd_sc_hd__clkbuf_1 _18744_ (.A(_02932_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _18745_ (.A0(_01362_),
    .A1(\core.decoded_imm_j[19] ),
    .S(_04978_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _18746_ (.A(_02933_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _18747_ (.A0(net25),
    .A1(_10238_),
    .S(_02913_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _18748_ (.A(_02934_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _18749_ (.A0(_01374_),
    .A1(_07200_),
    .S(_02925_),
    .X(_02935_));
 sky130_fd_sc_hd__buf_1 _18750_ (.A(_02935_),
    .X(_00761_));
 sky130_fd_sc_hd__inv_2 _18751_ (.A(_01349_),
    .Y(_02936_));
 sky130_fd_sc_hd__and4_1 _18752_ (.A(_10023_),
    .B(_10013_),
    .C(_02936_),
    .D(_10010_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(_02937_),
    .A1(\core.is_lb_lh_lw_lbu_lhu ),
    .S(_02925_),
    .X(_02938_));
 sky130_fd_sc_hd__buf_2 _18754_ (.A(_02938_),
    .X(_00762_));
 sky130_fd_sc_hd__a2bb2o_1 _18755_ (.A1_N(_10058_),
    .A2_N(_10245_),
    .B1(_10249_),
    .B2(_10268_),
    .X(_02939_));
 sky130_fd_sc_hd__inv_2 _18756_ (.A(_10221_),
    .Y(_02940_));
 sky130_fd_sc_hd__a22o_1 _18757_ (.A1(_04519_),
    .A2(_10218_),
    .B1(_02939_),
    .B2(_02940_),
    .X(_00763_));
 sky130_fd_sc_hd__nand2_1 _18758_ (.A(_10247_),
    .B(_04425_),
    .Y(_02941_));
 sky130_fd_sc_hd__and2_1 _18759_ (.A(_10058_),
    .B(\core.is_alu_reg_imm ),
    .X(_02942_));
 sky130_fd_sc_hd__o22a_1 _18760_ (.A1(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .A2(_10247_),
    .B1(_02941_),
    .B2(_02942_),
    .X(_00764_));
 sky130_fd_sc_hd__and4_1 _18761_ (.A(_10023_),
    .B(_01348_),
    .C(_02936_),
    .D(_10010_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _18762_ (.A0(_02943_),
    .A1(_04468_),
    .S(_02925_),
    .X(_02944_));
 sky130_fd_sc_hd__buf_1 _18763_ (.A(_02944_),
    .X(_00765_));
 sky130_fd_sc_hd__nor2_1 _18764_ (.A(_04477_),
    .B(_10247_),
    .Y(_02945_));
 sky130_fd_sc_hd__a31o_1 _18765_ (.A1(_02939_),
    .A2(\core.is_alu_reg_reg ),
    .A3(_10247_),
    .B1(_02945_),
    .X(_00766_));
 sky130_fd_sc_hd__or3b_1 _18766_ (.A(_10024_),
    .B(_04978_),
    .C_N(_10150_),
    .X(_02946_));
 sky130_fd_sc_hd__nand2_1 _18767_ (.A(_04979_),
    .B(_04975_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21oi_1 _18768_ (.A1(_02946_),
    .A2(_02947_),
    .B1(_10256_),
    .Y(_00767_));
 sky130_fd_sc_hd__clkbuf_2 _18769_ (.A(_04364_),
    .X(_02948_));
 sky130_fd_sc_hd__or3_1 _18770_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .B(\core.is_sb_sh_sw ),
    .C(_02900_),
    .X(_02949_));
 sky130_fd_sc_hd__nand2_1 _18771_ (.A(_02949_),
    .B(_10238_),
    .Y(_02950_));
 sky130_fd_sc_hd__o21a_1 _18772_ (.A1(_06657_),
    .A2(_07202_),
    .B1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__buf_1 _18773_ (.A(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_2 _18774_ (.A(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o21ai_4 _18775_ (.A1(_10265_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__mux2_1 _18776_ (.A0(_02954_),
    .A1(\core.decoded_imm[31] ),
    .S(_02903_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _18777_ (.A(_02955_),
    .X(_00768_));
 sky130_fd_sc_hd__o21ai_1 _18778_ (.A1(_10266_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02956_));
 sky130_fd_sc_hd__mux2_1 _18779_ (.A0(_02956_),
    .A1(\core.decoded_imm[30] ),
    .S(_02903_),
    .X(_02957_));
 sky130_fd_sc_hd__buf_1 _18780_ (.A(_02957_),
    .X(_00769_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18781_ (.A(_04365_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_4 _18782_ (.A(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__a21bo_1 _18783_ (.A1(\core.mem_rdata_q[29] ),
    .A2(_02959_),
    .B1_N(_02952_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _18784_ (.A0(_02960_),
    .A1(\core.decoded_imm[29] ),
    .S(_02903_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _18785_ (.A(_02961_),
    .X(_00770_));
 sky130_fd_sc_hd__o21ai_1 _18786_ (.A1(_10241_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02962_));
 sky130_fd_sc_hd__mux2_1 _18787_ (.A0(_02962_),
    .A1(\core.decoded_imm[28] ),
    .S(_02903_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_1 _18788_ (.A(_02963_),
    .X(_00771_));
 sky130_fd_sc_hd__o21ai_1 _18789_ (.A1(_10294_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02964_));
 sky130_fd_sc_hd__mux2_1 _18790_ (.A0(_02964_),
    .A1(\core.decoded_imm[27] ),
    .S(_02903_),
    .X(_02965_));
 sky130_fd_sc_hd__buf_1 _18791_ (.A(_02965_),
    .X(_00772_));
 sky130_fd_sc_hd__a21bo_1 _18792_ (.A1(\core.mem_rdata_q[26] ),
    .A2(_02959_),
    .B1_N(_02952_),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_4 _18793_ (.A(_10215_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _18794_ (.A0(_02966_),
    .A1(\core.decoded_imm[26] ),
    .S(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_2 _18795_ (.A(_02968_),
    .X(_00773_));
 sky130_fd_sc_hd__o21ai_2 _18796_ (.A1(_10240_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02969_));
 sky130_fd_sc_hd__mux2_1 _18797_ (.A0(_02969_),
    .A1(\core.decoded_imm[25] ),
    .S(_02967_),
    .X(_02970_));
 sky130_fd_sc_hd__buf_1 _18798_ (.A(_02970_),
    .X(_00774_));
 sky130_fd_sc_hd__o21ai_1 _18799_ (.A1(_10293_),
    .A2(_02948_),
    .B1(_02953_),
    .Y(_02971_));
 sky130_fd_sc_hd__mux2_1 _18800_ (.A0(_02971_),
    .A1(\core.decoded_imm[24] ),
    .S(_02967_),
    .X(_02972_));
 sky130_fd_sc_hd__buf_1 _18801_ (.A(_02972_),
    .X(_00775_));
 sky130_fd_sc_hd__o21ai_1 _18802_ (.A1(_10304_),
    .A2(_04364_),
    .B1(_02952_),
    .Y(_02973_));
 sky130_fd_sc_hd__mux2_1 _18803_ (.A0(_02973_),
    .A1(\core.decoded_imm[23] ),
    .S(_02967_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _18804_ (.A(_02974_),
    .X(_00776_));
 sky130_fd_sc_hd__o21ai_1 _18805_ (.A1(_10303_),
    .A2(_04364_),
    .B1(_02952_),
    .Y(_02975_));
 sky130_fd_sc_hd__mux2_1 _18806_ (.A0(_02975_),
    .A1(\core.decoded_imm[22] ),
    .S(_02967_),
    .X(_02976_));
 sky130_fd_sc_hd__clkbuf_1 _18807_ (.A(_02976_),
    .X(_00777_));
 sky130_fd_sc_hd__o21ai_1 _18808_ (.A1(_10302_),
    .A2(_04364_),
    .B1(_02952_),
    .Y(_02977_));
 sky130_fd_sc_hd__mux2_1 _18809_ (.A0(_02977_),
    .A1(\core.decoded_imm[21] ),
    .S(_02967_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_1 _18810_ (.A(_02978_),
    .X(_00778_));
 sky130_fd_sc_hd__a21bo_1 _18811_ (.A1(\core.mem_rdata_q[20] ),
    .A2(_02959_),
    .B1_N(_02951_),
    .X(_02979_));
 sky130_fd_sc_hd__buf_2 _18812_ (.A(_10215_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _18813_ (.A0(_02979_),
    .A1(\core.decoded_imm[20] ),
    .S(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _18814_ (.A(_02981_),
    .X(_00779_));
 sky130_fd_sc_hd__inv_2 _18815_ (.A(_02950_),
    .Y(_02982_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18816_ (.A(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__a221o_1 _18817_ (.A1(_06949_),
    .A2(\core.decoded_imm_j[19] ),
    .B1(\core.mem_rdata_q[19] ),
    .B2(_02959_),
    .C1(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _18818_ (.A0(_02984_),
    .A1(\core.decoded_imm[19] ),
    .S(_02980_),
    .X(_02985_));
 sky130_fd_sc_hd__buf_1 _18819_ (.A(_02985_),
    .X(_00780_));
 sky130_fd_sc_hd__a221o_1 _18820_ (.A1(_06949_),
    .A2(\core.decoded_imm_j[18] ),
    .B1(\core.mem_rdata_q[18] ),
    .B2(_02959_),
    .C1(_02983_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _18821_ (.A0(_02986_),
    .A1(\core.decoded_imm[18] ),
    .S(_02980_),
    .X(_02987_));
 sky130_fd_sc_hd__clkbuf_1 _18822_ (.A(_02987_),
    .X(_00781_));
 sky130_fd_sc_hd__a221o_1 _18823_ (.A1(_06949_),
    .A2(\core.decoded_imm_j[17] ),
    .B1(\core.mem_rdata_q[17] ),
    .B2(_02959_),
    .C1(_02983_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _18824_ (.A0(_02988_),
    .A1(\core.decoded_imm[17] ),
    .S(_02980_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _18825_ (.A(_02989_),
    .X(_00782_));
 sky130_fd_sc_hd__a221o_1 _18826_ (.A1(_06949_),
    .A2(\core.decoded_imm_j[16] ),
    .B1(\core.mem_rdata_q[16] ),
    .B2(_02958_),
    .C1(_02983_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _18827_ (.A0(_02990_),
    .A1(\core.decoded_imm[16] ),
    .S(_02980_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _18828_ (.A(_02991_),
    .X(_00783_));
 sky130_fd_sc_hd__a221o_1 _18829_ (.A1(_06949_),
    .A2(\core.decoded_imm_j[15] ),
    .B1(\core.mem_rdata_q[15] ),
    .B2(_02958_),
    .C1(_02983_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _18830_ (.A0(_02992_),
    .A1(\core.decoded_imm[15] ),
    .S(_02980_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _18831_ (.A(_02993_),
    .X(_00784_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18832_ (.A(_06607_),
    .X(_02994_));
 sky130_fd_sc_hd__a221o_1 _18833_ (.A1(_02994_),
    .A2(\core.decoded_imm_j[14] ),
    .B1(\core.mem_rdata_q[14] ),
    .B2(_02958_),
    .C1(_02983_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_2 _18834_ (.A(_10215_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _18835_ (.A0(_02995_),
    .A1(\core.decoded_imm[14] ),
    .S(_02996_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _18836_ (.A(_02997_),
    .X(_00785_));
 sky130_fd_sc_hd__a221o_1 _18837_ (.A1(_02994_),
    .A2(\core.decoded_imm_j[13] ),
    .B1(\core.mem_rdata_q[13] ),
    .B2(_02958_),
    .C1(_02982_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_8 _18838_ (.A0(_02998_),
    .A1(\core.decoded_imm[13] ),
    .S(_02996_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _18839_ (.A(_02999_),
    .X(_00786_));
 sky130_fd_sc_hd__a221o_1 _18840_ (.A1(_02994_),
    .A2(\core.decoded_imm_j[12] ),
    .B1(\core.mem_rdata_q[12] ),
    .B2(_02958_),
    .C1(_02982_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _18841_ (.A0(_03000_),
    .A1(\core.decoded_imm[12] ),
    .S(_02996_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _18842_ (.A(_03001_),
    .X(_00787_));
 sky130_fd_sc_hd__a22o_1 _18843_ (.A1(_06607_),
    .A2(_04577_),
    .B1(_04467_),
    .B2(_10238_),
    .X(_03002_));
 sky130_fd_sc_hd__a221o_1 _18844_ (.A1(_04975_),
    .A2(\core.mem_rdata_q[7] ),
    .B1(_02901_),
    .B2(_10238_),
    .C1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _18845_ (.A0(_03003_),
    .A1(\core.decoded_imm[11] ),
    .S(_02996_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _18846_ (.A(_03004_),
    .X(_00788_));
 sky130_fd_sc_hd__clkbuf_4 _18847_ (.A(_02949_),
    .X(_03005_));
 sky130_fd_sc_hd__a22o_1 _18848_ (.A1(_06973_),
    .A2(\core.decoded_imm_j[10] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[30] ),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _18849_ (.A0(_03006_),
    .A1(\core.decoded_imm[10] ),
    .S(_02996_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _18850_ (.A(_03007_),
    .X(_00789_));
 sky130_fd_sc_hd__a22o_1 _18851_ (.A1(_06973_),
    .A2(\core.decoded_imm_j[9] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[29] ),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _18852_ (.A0(_03008_),
    .A1(\core.decoded_imm[9] ),
    .S(_02996_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _18853_ (.A(_03009_),
    .X(_00790_));
 sky130_fd_sc_hd__a22o_1 _18854_ (.A1(_06897_),
    .A2(\core.decoded_imm_j[8] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[28] ),
    .X(_03010_));
 sky130_fd_sc_hd__buf_2 _18855_ (.A(_10215_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _18856_ (.A0(_03010_),
    .A1(\core.decoded_imm[8] ),
    .S(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _18857_ (.A(_03012_),
    .X(_00791_));
 sky130_fd_sc_hd__a22o_1 _18858_ (.A1(_06897_),
    .A2(\core.decoded_imm_j[7] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[27] ),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _18859_ (.A0(_03013_),
    .A1(\core.decoded_imm[7] ),
    .S(_03011_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _18860_ (.A(_03014_),
    .X(_00792_));
 sky130_fd_sc_hd__a22o_1 _18861_ (.A1(_06897_),
    .A2(\core.decoded_imm_j[6] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[26] ),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _18862_ (.A0(_03015_),
    .A1(\core.decoded_imm[6] ),
    .S(_03011_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _18863_ (.A(_03016_),
    .X(_00793_));
 sky130_fd_sc_hd__a22o_1 _18864_ (.A1(_06897_),
    .A2(\core.decoded_imm_j[5] ),
    .B1(_03005_),
    .B2(\core.mem_rdata_q[25] ),
    .X(_03017_));
 sky130_fd_sc_hd__mux2_1 _18865_ (.A0(_03017_),
    .A1(\core.decoded_imm[5] ),
    .S(_03011_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _18866_ (.A(_03018_),
    .X(_00794_));
 sky130_fd_sc_hd__o21a_1 _18867_ (.A1(_04488_),
    .A2(_04467_),
    .B1(\core.mem_rdata_q[11] ),
    .X(_03019_));
 sky130_fd_sc_hd__a221o_1 _18868_ (.A1(_02994_),
    .A2(_04576_),
    .B1(_02901_),
    .B2(\core.mem_rdata_q[24] ),
    .C1(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _18869_ (.A0(_03020_),
    .A1(\core.decoded_imm[4] ),
    .S(_03011_),
    .X(_03021_));
 sky130_fd_sc_hd__buf_1 _18870_ (.A(_03021_),
    .X(_00795_));
 sky130_fd_sc_hd__o21a_1 _18871_ (.A1(_04488_),
    .A2(_04467_),
    .B1(\core.mem_rdata_q[10] ),
    .X(_03022_));
 sky130_fd_sc_hd__a221o_1 _18872_ (.A1(_02994_),
    .A2(_04575_),
    .B1(_02901_),
    .B2(\core.mem_rdata_q[23] ),
    .C1(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _18873_ (.A0(_03023_),
    .A1(\core.decoded_imm[3] ),
    .S(_03011_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _18874_ (.A(_03024_),
    .X(_00796_));
 sky130_fd_sc_hd__o21a_1 _18875_ (.A1(_04488_),
    .A2(_04467_),
    .B1(\core.mem_rdata_q[9] ),
    .X(_03025_));
 sky130_fd_sc_hd__a221o_1 _18876_ (.A1(_02994_),
    .A2(\core.decoded_imm_j[2] ),
    .B1(_02901_),
    .B2(\core.mem_rdata_q[22] ),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _18877_ (.A0(_03026_),
    .A1(\core.decoded_imm[2] ),
    .S(_10226_),
    .X(_03027_));
 sky130_fd_sc_hd__buf_1 _18878_ (.A(_03027_),
    .X(_00797_));
 sky130_fd_sc_hd__o21a_1 _18879_ (.A1(_04488_),
    .A2(_04467_),
    .B1(\core.mem_rdata_q[8] ),
    .X(_03028_));
 sky130_fd_sc_hd__a221o_1 _18880_ (.A1(_06703_),
    .A2(_05942_),
    .B1(_02901_),
    .B2(\core.mem_rdata_q[21] ),
    .C1(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _18881_ (.A0(_03029_),
    .A1(\core.decoded_imm[1] ),
    .S(_10226_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _18882_ (.A(_03030_),
    .X(_00798_));
 sky130_fd_sc_hd__or3_1 _18883_ (.A(\core.latched_rd[3] ),
    .B(\core.latched_rd[2] ),
    .C(_09317_),
    .X(_03031_));
 sky130_fd_sc_hd__nor2_1 _18884_ (.A(_03031_),
    .B(_02778_),
    .Y(_03032_));
 sky130_fd_sc_hd__buf_4 _18885_ (.A(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_2 _18886_ (.A(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_2 _18887_ (.A0(\core.cpuregs[17][0] ),
    .A1(_10062_),
    .S(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _18888_ (.A(_03035_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_4 _18889_ (.A0(\core.cpuregs[17][1] ),
    .A1(_10069_),
    .S(_03034_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_2 _18890_ (.A(_03036_),
    .X(_00800_));
 sky130_fd_sc_hd__buf_2 _18891_ (.A(_03033_),
    .X(_03037_));
 sky130_fd_sc_hd__mux2_1 _18892_ (.A0(\core.cpuregs[17][2] ),
    .A1(_10071_),
    .S(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _18893_ (.A(_03038_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _18894_ (.A0(\core.cpuregs[17][3] ),
    .A1(_10074_),
    .S(_03037_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_1 _18895_ (.A(_03039_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _18896_ (.A0(\core.cpuregs[17][4] ),
    .A1(_10076_),
    .S(_03037_),
    .X(_03040_));
 sky130_fd_sc_hd__buf_1 _18897_ (.A(_03040_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _18898_ (.A0(\core.cpuregs[17][5] ),
    .A1(_10078_),
    .S(_03037_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _18899_ (.A(_03041_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _18900_ (.A0(\core.cpuregs[17][6] ),
    .A1(_10080_),
    .S(_03037_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _18901_ (.A(_03042_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _18902_ (.A0(\core.cpuregs[17][7] ),
    .A1(_10082_),
    .S(_03037_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _18903_ (.A(_03043_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _18904_ (.A0(\core.cpuregs[17][8] ),
    .A1(_10084_),
    .S(_03033_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_2 _18905_ (.A(_03044_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _18906_ (.A0(\core.cpuregs[17][9] ),
    .A1(_10086_),
    .S(_03033_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _18907_ (.A(_03045_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _18908_ (.A0(\core.cpuregs[17][10] ),
    .A1(_10088_),
    .S(_03033_),
    .X(_03046_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _18909_ (.A(_03046_),
    .X(_00809_));
 sky130_fd_sc_hd__inv_2 _18910_ (.A(_03032_),
    .Y(_03047_));
 sky130_fd_sc_hd__clkbuf_2 _18911_ (.A(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _18912_ (.A0(_10090_),
    .A1(\core.cpuregs[17][11] ),
    .S(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _18913_ (.A(_03049_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _18914_ (.A0(\core.cpuregs[17][12] ),
    .A1(_10094_),
    .S(_03033_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_1 _18915_ (.A(_03050_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _18916_ (.A0(_10096_),
    .A1(\core.cpuregs[17][13] ),
    .S(_03048_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _18917_ (.A(_03051_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _18918_ (.A0(_10098_),
    .A1(\core.cpuregs[17][14] ),
    .S(_03047_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _18919_ (.A(_03052_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(_10100_),
    .A1(\core.cpuregs[17][15] ),
    .S(_03047_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _18921_ (.A(_03053_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_2 _18922_ (.A0(_10102_),
    .A1(\core.cpuregs[17][16] ),
    .S(_03047_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _18923_ (.A(_03054_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(_10104_),
    .A1(\core.cpuregs[17][17] ),
    .S(_03047_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_2 _18925_ (.A(_03055_),
    .X(_00816_));
 sky130_fd_sc_hd__and2_1 _18926_ (.A(_03048_),
    .B(\core.cpuregs[17][18] ),
    .X(_03056_));
 sky130_fd_sc_hd__a21o_1 _18927_ (.A1(_09779_),
    .A2(_03034_),
    .B1(_03056_),
    .X(_00817_));
 sky130_fd_sc_hd__clkbuf_4 _18928_ (.A(_03034_),
    .X(_03057_));
 sky130_fd_sc_hd__nand2_2 _18929_ (.A(_10107_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__clkbuf_2 _18930_ (.A(_03048_),
    .X(_03059_));
 sky130_fd_sc_hd__nand2_1 _18931_ (.A(_03059_),
    .B(net127),
    .Y(_03060_));
 sky130_fd_sc_hd__nand2_1 _18932_ (.A(_03058_),
    .B(_03060_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _18933_ (.A(_10112_),
    .B(_03057_),
    .Y(_03061_));
 sky130_fd_sc_hd__nand2_1 _18934_ (.A(_03059_),
    .B(\core.cpuregs[17][20] ),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_1 _18935_ (.A(_03061_),
    .B(_03062_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _18936_ (.A(_10115_),
    .B(_03057_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _18937_ (.A(_03059_),
    .B(net120),
    .Y(_03064_));
 sky130_fd_sc_hd__nand2_1 _18938_ (.A(_03063_),
    .B(_03064_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_1 _18939_ (.A(_10118_),
    .B(_03057_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _18940_ (.A(_03059_),
    .B(\core.cpuregs[17][22] ),
    .Y(_03066_));
 sky130_fd_sc_hd__nand2_1 _18941_ (.A(_03065_),
    .B(_03066_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _18942_ (.A(_10121_),
    .B(_03057_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_4 _18943_ (.A(_03059_),
    .B(\core.cpuregs[17][23] ),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_1 _18944_ (.A(_03067_),
    .B(_03068_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_1 _18945_ (.A(_10124_),
    .B(_03057_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_1 _18946_ (.A(_03059_),
    .B(\core.cpuregs[17][24] ),
    .Y(_03070_));
 sky130_fd_sc_hd__nand2_1 _18947_ (.A(_03069_),
    .B(_03070_),
    .Y(_00823_));
 sky130_fd_sc_hd__clkbuf_2 _18948_ (.A(_03034_),
    .X(_03071_));
 sky130_fd_sc_hd__nand2_4 _18949_ (.A(_10127_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__clkbuf_4 _18950_ (.A(_03048_),
    .X(_03073_));
 sky130_fd_sc_hd__nand2_4 _18951_ (.A(_03073_),
    .B(\core.cpuregs[17][25] ),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _18952_ (.A(_03072_),
    .B(_03074_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _18953_ (.A(_10132_),
    .B(_03071_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_1 _18954_ (.A(_03073_),
    .B(\core.cpuregs[17][26] ),
    .Y(_03076_));
 sky130_fd_sc_hd__nand2_1 _18955_ (.A(_03075_),
    .B(_03076_),
    .Y(_00825_));
 sky130_fd_sc_hd__nand2_1 _18956_ (.A(_10135_),
    .B(_03071_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2_1 _18957_ (.A(_03073_),
    .B(\core.cpuregs[17][27] ),
    .Y(_03078_));
 sky130_fd_sc_hd__nand2_1 _18958_ (.A(_03077_),
    .B(_03078_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _18959_ (.A(_10138_),
    .B(_03071_),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_4 _18960_ (.A(_03073_),
    .B(\core.cpuregs[17][28] ),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2_1 _18961_ (.A(_03079_),
    .B(_03080_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_2 _18962_ (.A(_10141_),
    .B(_03071_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand2_4 _18963_ (.A(_03073_),
    .B(\core.cpuregs[17][29] ),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _18964_ (.A(_03081_),
    .B(_03082_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _18965_ (.A(_10144_),
    .B(_03071_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_4 _18966_ (.A(_03073_),
    .B(\core.cpuregs[17][30] ),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _18967_ (.A(_03083_),
    .B(_03084_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_1 _18968_ (.A(_10147_),
    .B(_03034_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _18969_ (.A(_03048_),
    .B(\core.cpuregs[17][31] ),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _18970_ (.A(_03085_),
    .B(_03086_),
    .Y(_00830_));
 sky130_fd_sc_hd__clkbuf_2 _18971_ (.A(_09314_),
    .X(_03087_));
 sky130_fd_sc_hd__nor2_1 _18972_ (.A(_03031_),
    .B(_09950_),
    .Y(_03088_));
 sky130_fd_sc_hd__clkbuf_2 _18973_ (.A(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_2 _18974_ (.A(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _18975_ (.A0(\core.cpuregs[16][0] ),
    .A1(_03087_),
    .S(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_8 _18976_ (.A(_03091_),
    .X(_00831_));
 sky130_fd_sc_hd__buf_1 _18977_ (.A(_09336_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _18978_ (.A0(\core.cpuregs[16][1] ),
    .A1(_03092_),
    .S(_03090_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _18979_ (.A(_03093_),
    .X(_00832_));
 sky130_fd_sc_hd__buf_1 _18980_ (.A(_09339_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_4 _18981_ (.A(_03089_),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _18982_ (.A0(\core.cpuregs[16][2] ),
    .A1(_03094_),
    .S(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _18983_ (.A(_03096_),
    .X(_00833_));
 sky130_fd_sc_hd__buf_2 _18984_ (.A(_09348_),
    .X(_03097_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(\core.cpuregs[16][3] ),
    .A1(_03097_),
    .S(_03095_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _18986_ (.A(_03098_),
    .X(_00834_));
 sky130_fd_sc_hd__buf_2 _18987_ (.A(_09356_),
    .X(_03099_));
 sky130_fd_sc_hd__mux2_1 _18988_ (.A0(\core.cpuregs[16][4] ),
    .A1(_03099_),
    .S(_03095_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _18989_ (.A(_03100_),
    .X(_00835_));
 sky130_fd_sc_hd__clkbuf_2 _18990_ (.A(_09362_),
    .X(_03101_));
 sky130_fd_sc_hd__mux2_1 _18991_ (.A0(\core.cpuregs[16][5] ),
    .A1(_03101_),
    .S(_03095_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _18992_ (.A(_03102_),
    .X(_00836_));
 sky130_fd_sc_hd__buf_2 _18993_ (.A(_09368_),
    .X(_03103_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(\core.cpuregs[16][6] ),
    .A1(_03103_),
    .S(_03095_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _18995_ (.A(_03104_),
    .X(_00837_));
 sky130_fd_sc_hd__buf_2 _18996_ (.A(_09374_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _18997_ (.A0(\core.cpuregs[16][7] ),
    .A1(_03105_),
    .S(_03095_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _18998_ (.A(_03106_),
    .X(_00838_));
 sky130_fd_sc_hd__clkbuf_4 _18999_ (.A(_09380_),
    .X(_03107_));
 sky130_fd_sc_hd__mux2_1 _19000_ (.A0(\core.cpuregs[16][8] ),
    .A1(_03107_),
    .S(_03089_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_2 _19001_ (.A(_03108_),
    .X(_00839_));
 sky130_fd_sc_hd__buf_4 _19002_ (.A(_09387_),
    .X(_03109_));
 sky130_fd_sc_hd__mux2_1 _19003_ (.A0(\core.cpuregs[16][9] ),
    .A1(_03109_),
    .S(_03089_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_1 _19004_ (.A(_03110_),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_4 _19005_ (.A(_09394_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _19006_ (.A0(\core.cpuregs[16][10] ),
    .A1(_03111_),
    .S(_03089_),
    .X(_03112_));
 sky130_fd_sc_hd__clkbuf_1 _19007_ (.A(_03112_),
    .X(_00841_));
 sky130_fd_sc_hd__buf_1 _19008_ (.A(_09400_),
    .X(_03113_));
 sky130_fd_sc_hd__inv_2 _19009_ (.A(_03088_),
    .Y(_03114_));
 sky130_fd_sc_hd__buf_4 _19010_ (.A(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__mux2_1 _19011_ (.A0(_03113_),
    .A1(\core.cpuregs[16][11] ),
    .S(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__clkbuf_1 _19012_ (.A(_03116_),
    .X(_00842_));
 sky130_fd_sc_hd__buf_1 _19013_ (.A(_09407_),
    .X(_03117_));
 sky130_fd_sc_hd__mux2_1 _19014_ (.A0(\core.cpuregs[16][12] ),
    .A1(_03117_),
    .S(_03089_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _19015_ (.A(_03118_),
    .X(_00843_));
 sky130_fd_sc_hd__buf_2 _19016_ (.A(_09413_),
    .X(_03119_));
 sky130_fd_sc_hd__mux2_1 _19017_ (.A0(_03119_),
    .A1(\core.cpuregs[16][13] ),
    .S(_03115_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_2 _19018_ (.A(_03120_),
    .X(_00844_));
 sky130_fd_sc_hd__buf_1 _19019_ (.A(_09418_),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_2 _19020_ (.A0(_03121_),
    .A1(\core.cpuregs[16][14] ),
    .S(_03114_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _19021_ (.A(_03122_),
    .X(_00845_));
 sky130_fd_sc_hd__buf_2 _19022_ (.A(_09423_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _19023_ (.A0(_03123_),
    .A1(\core.cpuregs[16][15] ),
    .S(_03114_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _19024_ (.A(_03124_),
    .X(_00846_));
 sky130_fd_sc_hd__buf_2 _19025_ (.A(_09430_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _19026_ (.A0(_03125_),
    .A1(\core.cpuregs[16][16] ),
    .S(_03114_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _19027_ (.A(_03126_),
    .X(_00847_));
 sky130_fd_sc_hd__buf_2 _19028_ (.A(_09435_),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_1 _19029_ (.A0(_03127_),
    .A1(\core.cpuregs[16][17] ),
    .S(_03114_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _19030_ (.A(_03128_),
    .X(_00848_));
 sky130_fd_sc_hd__and2_1 _19031_ (.A(_03115_),
    .B(\core.cpuregs[16][18] ),
    .X(_03129_));
 sky130_fd_sc_hd__a21o_1 _19032_ (.A1(_09779_),
    .A2(_03090_),
    .B1(_03129_),
    .X(_00849_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19033_ (.A(_09447_),
    .X(_03130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19034_ (.A(_03090_),
    .X(_03131_));
 sky130_fd_sc_hd__nand2_1 _19035_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19036_ (.A(_03115_),
    .X(_03133_));
 sky130_fd_sc_hd__nand2_2 _19037_ (.A(_03133_),
    .B(\core.cpuregs[16][19] ),
    .Y(_03134_));
 sky130_fd_sc_hd__nand2_1 _19038_ (.A(_03132_),
    .B(_03134_),
    .Y(_00850_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19039_ (.A(_09457_),
    .X(_03135_));
 sky130_fd_sc_hd__nand2_1 _19040_ (.A(_03135_),
    .B(_03131_),
    .Y(_03136_));
 sky130_fd_sc_hd__nand2_1 _19041_ (.A(_03133_),
    .B(\core.cpuregs[16][20] ),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _19042_ (.A(_03136_),
    .B(_03137_),
    .Y(_00851_));
 sky130_fd_sc_hd__clkbuf_2 _19043_ (.A(_09466_),
    .X(_03138_));
 sky130_fd_sc_hd__nand2_1 _19044_ (.A(_03138_),
    .B(_03131_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _19045_ (.A(_03133_),
    .B(\core.cpuregs[16][21] ),
    .Y(_03140_));
 sky130_fd_sc_hd__nand2_1 _19046_ (.A(_03139_),
    .B(_03140_),
    .Y(_00852_));
 sky130_fd_sc_hd__clkbuf_4 _19047_ (.A(_09473_),
    .X(_03141_));
 sky130_fd_sc_hd__nand2_2 _19048_ (.A(_03141_),
    .B(_03131_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _19049_ (.A(_03133_),
    .B(\core.cpuregs[16][22] ),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _19050_ (.A(_03142_),
    .B(_03143_),
    .Y(_00853_));
 sky130_fd_sc_hd__buf_6 _19051_ (.A(_09480_),
    .X(_03144_));
 sky130_fd_sc_hd__nand2_1 _19052_ (.A(_03144_),
    .B(_03131_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _19053_ (.A(_03133_),
    .B(\core.cpuregs[16][23] ),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _19054_ (.A(_03145_),
    .B(_03146_),
    .Y(_00854_));
 sky130_fd_sc_hd__buf_6 _19055_ (.A(_09488_),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_1 _19056_ (.A(_03147_),
    .B(_03131_),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_1 _19057_ (.A(_03133_),
    .B(\core.cpuregs[16][24] ),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _19058_ (.A(_03148_),
    .B(_03149_),
    .Y(_00855_));
 sky130_fd_sc_hd__clkbuf_2 _19059_ (.A(_09498_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_2 _19060_ (.A(_03090_),
    .X(_03151_));
 sky130_fd_sc_hd__nand2_1 _19061_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19062_ (.A(_03115_),
    .X(_03153_));
 sky130_fd_sc_hd__nand2_1 _19063_ (.A(_03153_),
    .B(\core.cpuregs[16][25] ),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _19064_ (.A(_03152_),
    .B(_03154_),
    .Y(_00856_));
 sky130_fd_sc_hd__clkbuf_4 _19065_ (.A(_09508_),
    .X(_03155_));
 sky130_fd_sc_hd__nand2_2 _19066_ (.A(_03155_),
    .B(_03151_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand2_1 _19067_ (.A(_03153_),
    .B(\core.cpuregs[16][26] ),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _19068_ (.A(_03156_),
    .B(_03157_),
    .Y(_00857_));
 sky130_fd_sc_hd__buf_2 _19069_ (.A(_09515_),
    .X(_03158_));
 sky130_fd_sc_hd__nand2_1 _19070_ (.A(_03158_),
    .B(_03151_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _19071_ (.A(_03153_),
    .B(\core.cpuregs[16][27] ),
    .Y(_03160_));
 sky130_fd_sc_hd__nand2_1 _19072_ (.A(_03159_),
    .B(_03160_),
    .Y(_00858_));
 sky130_fd_sc_hd__buf_6 _19073_ (.A(_09524_),
    .X(_03161_));
 sky130_fd_sc_hd__nand2_1 _19074_ (.A(_03161_),
    .B(_03151_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_2 _19075_ (.A(_03153_),
    .B(\core.cpuregs[16][28] ),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_1 _19076_ (.A(_03162_),
    .B(_03163_),
    .Y(_00859_));
 sky130_fd_sc_hd__clkbuf_2 _19077_ (.A(_09533_),
    .X(_03164_));
 sky130_fd_sc_hd__nand2_1 _19078_ (.A(_03164_),
    .B(_03151_),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_1 _19079_ (.A(_03153_),
    .B(\core.cpuregs[16][29] ),
    .Y(_03166_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(_03165_),
    .B(_03166_),
    .Y(_00860_));
 sky130_fd_sc_hd__buf_6 _19081_ (.A(_09541_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_1 _19082_ (.A(_03167_),
    .B(_03151_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_1 _19083_ (.A(_03153_),
    .B(\core.cpuregs[16][30] ),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _19084_ (.A(_03168_),
    .B(_03169_),
    .Y(_00861_));
 sky130_fd_sc_hd__clkbuf_2 _19085_ (.A(_09550_),
    .X(_03170_));
 sky130_fd_sc_hd__nand2_1 _19086_ (.A(_03170_),
    .B(_03090_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _19087_ (.A(_03115_),
    .B(\core.cpuregs[16][31] ),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_1 _19088_ (.A(_03171_),
    .B(_03172_),
    .Y(_00862_));
 sky130_fd_sc_hd__or3_4 _19089_ (.A(\core.latched_rd[4] ),
    .B(_09318_),
    .C(_09319_),
    .X(_03173_));
 sky130_fd_sc_hd__nor2_1 _19090_ (.A(_03173_),
    .B(_09812_),
    .Y(_03174_));
 sky130_fd_sc_hd__clkbuf_4 _19091_ (.A(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_2 _19092_ (.A(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__mux2_1 _19093_ (.A0(\core.cpuregs[15][0] ),
    .A1(_03087_),
    .S(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__buf_1 _19094_ (.A(_03177_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _19095_ (.A0(\core.cpuregs[15][1] ),
    .A1(_03092_),
    .S(_03176_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _19096_ (.A(_03178_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_2 _19097_ (.A(_03175_),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_2 _19098_ (.A0(\core.cpuregs[15][2] ),
    .A1(_03094_),
    .S(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _19099_ (.A(_03180_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _19100_ (.A0(\core.cpuregs[15][3] ),
    .A1(_03097_),
    .S(_03179_),
    .X(_03181_));
 sky130_fd_sc_hd__buf_2 _19101_ (.A(_03181_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _19102_ (.A0(\core.cpuregs[15][4] ),
    .A1(_03099_),
    .S(_03179_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _19103_ (.A(_03182_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _19104_ (.A0(\core.cpuregs[15][5] ),
    .A1(_03101_),
    .S(_03179_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_4 _19105_ (.A(_03183_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _19106_ (.A0(\core.cpuregs[15][6] ),
    .A1(_03103_),
    .S(_03179_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _19107_ (.A(_03184_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _19108_ (.A0(\core.cpuregs[15][7] ),
    .A1(_03105_),
    .S(_03179_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _19109_ (.A(_03185_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _19110_ (.A0(\core.cpuregs[15][8] ),
    .A1(_03107_),
    .S(_03175_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _19111_ (.A(_03186_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_2 _19112_ (.A0(\core.cpuregs[15][9] ),
    .A1(_03109_),
    .S(_03175_),
    .X(_03187_));
 sky130_fd_sc_hd__clkbuf_1 _19113_ (.A(_03187_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _19114_ (.A0(\core.cpuregs[15][10] ),
    .A1(_03111_),
    .S(_03175_),
    .X(_03188_));
 sky130_fd_sc_hd__clkbuf_1 _19115_ (.A(_03188_),
    .X(_00873_));
 sky130_fd_sc_hd__inv_2 _19116_ (.A(_03174_),
    .Y(_03189_));
 sky130_fd_sc_hd__clkbuf_4 _19117_ (.A(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _19118_ (.A0(_03113_),
    .A1(\core.cpuregs[15][11] ),
    .S(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__clkbuf_1 _19119_ (.A(_03191_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _19120_ (.A0(\core.cpuregs[15][12] ),
    .A1(_03117_),
    .S(_03175_),
    .X(_03192_));
 sky130_fd_sc_hd__clkbuf_1 _19121_ (.A(_03192_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _19122_ (.A0(_03119_),
    .A1(\core.cpuregs[15][13] ),
    .S(_03190_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_1 _19123_ (.A(_03193_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _19124_ (.A0(_03121_),
    .A1(\core.cpuregs[15][14] ),
    .S(_03189_),
    .X(_03194_));
 sky130_fd_sc_hd__clkbuf_1 _19125_ (.A(_03194_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _19126_ (.A0(_03123_),
    .A1(\core.cpuregs[15][15] ),
    .S(_03189_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _19127_ (.A(_03195_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _19128_ (.A0(_03125_),
    .A1(\core.cpuregs[15][16] ),
    .S(_03189_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_1 _19129_ (.A(_03196_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _19130_ (.A0(_03127_),
    .A1(\core.cpuregs[15][17] ),
    .S(_03189_),
    .X(_03197_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19131_ (.A(_03197_),
    .X(_00880_));
 sky130_fd_sc_hd__clkbuf_2 _19132_ (.A(_09441_),
    .X(_03198_));
 sky130_fd_sc_hd__nand2_1 _19133_ (.A(_03190_),
    .B(\core.cpuregs[15][18] ),
    .Y(_03199_));
 sky130_fd_sc_hd__a21bo_1 _19134_ (.A1(_03198_),
    .A2(_03176_),
    .B1_N(_03199_),
    .X(_00881_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19135_ (.A(_03176_),
    .X(_03200_));
 sky130_fd_sc_hd__nand2_1 _19136_ (.A(_03130_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__buf_2 _19137_ (.A(_03190_),
    .X(_03202_));
 sky130_fd_sc_hd__nand2_1 _19138_ (.A(_03202_),
    .B(net159),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _19139_ (.A(_03201_),
    .B(_03203_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _19140_ (.A(_03135_),
    .B(_03200_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand2_1 _19141_ (.A(_03202_),
    .B(\core.cpuregs[15][20] ),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _19142_ (.A(_03204_),
    .B(_03205_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _19143_ (.A(_03138_),
    .B(_03200_),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _19144_ (.A(_03202_),
    .B(net194),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _19145_ (.A(_03206_),
    .B(_03207_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _19146_ (.A(_03141_),
    .B(_03200_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _19147_ (.A(_03202_),
    .B(\core.cpuregs[15][22] ),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _19148_ (.A(_03208_),
    .B(_03209_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _19149_ (.A(_03144_),
    .B(_03200_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _19150_ (.A(_03202_),
    .B(\core.cpuregs[15][23] ),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_1 _19151_ (.A(_03210_),
    .B(_03211_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand2_1 _19152_ (.A(_03147_),
    .B(_03200_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _19153_ (.A(_03202_),
    .B(\core.cpuregs[15][24] ),
    .Y(_03213_));
 sky130_fd_sc_hd__nand2_1 _19154_ (.A(_03212_),
    .B(_03213_),
    .Y(_00887_));
 sky130_fd_sc_hd__clkbuf_4 _19155_ (.A(_03176_),
    .X(_03214_));
 sky130_fd_sc_hd__nand2_1 _19156_ (.A(_03150_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19157_ (.A(_03190_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _19158_ (.A(_03216_),
    .B(\core.cpuregs[15][25] ),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _19159_ (.A(_03215_),
    .B(_03217_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _19160_ (.A(_03155_),
    .B(_03214_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand2_1 _19161_ (.A(_03216_),
    .B(\core.cpuregs[15][26] ),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _19162_ (.A(_03218_),
    .B(_03219_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand2_1 _19163_ (.A(_03158_),
    .B(_03214_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_1 _19164_ (.A(_03216_),
    .B(\core.cpuregs[15][27] ),
    .Y(_03221_));
 sky130_fd_sc_hd__nand2_1 _19165_ (.A(_03220_),
    .B(_03221_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _19166_ (.A(_03161_),
    .B(_03214_),
    .Y(_03222_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(_03216_),
    .B(\core.cpuregs[15][28] ),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _19168_ (.A(_03222_),
    .B(_03223_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_2 _19169_ (.A(_03164_),
    .B(_03214_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _19170_ (.A(_03216_),
    .B(\core.cpuregs[15][29] ),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _19171_ (.A(_03224_),
    .B(_03225_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand2_1 _19172_ (.A(_03167_),
    .B(_03214_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _19173_ (.A(_03216_),
    .B(\core.cpuregs[15][30] ),
    .Y(_03227_));
 sky130_fd_sc_hd__nand2_1 _19174_ (.A(_03226_),
    .B(_03227_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand2_1 _19175_ (.A(_03170_),
    .B(_03176_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _19176_ (.A(_03190_),
    .B(\core.cpuregs[15][31] ),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _19177_ (.A(_03228_),
    .B(_03229_),
    .Y(_00894_));
 sky130_fd_sc_hd__nor2_1 _19178_ (.A(_03173_),
    .B(_10158_),
    .Y(_03230_));
 sky130_fd_sc_hd__clkbuf_4 _19179_ (.A(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_2 _19180_ (.A(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_2 _19181_ (.A0(\core.cpuregs[14][0] ),
    .A1(_03087_),
    .S(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__clkbuf_1 _19182_ (.A(_03233_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _19183_ (.A0(\core.cpuregs[14][1] ),
    .A1(_03092_),
    .S(_03232_),
    .X(_03234_));
 sky130_fd_sc_hd__clkbuf_1 _19184_ (.A(_03234_),
    .X(_00896_));
 sky130_fd_sc_hd__clkbuf_4 _19185_ (.A(_03231_),
    .X(_03235_));
 sky130_fd_sc_hd__mux2_1 _19186_ (.A0(\core.cpuregs[14][2] ),
    .A1(_03094_),
    .S(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_1 _19187_ (.A(_03236_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _19188_ (.A0(\core.cpuregs[14][3] ),
    .A1(_03097_),
    .S(_03235_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _19189_ (.A(_03237_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _19190_ (.A0(\core.cpuregs[14][4] ),
    .A1(_03099_),
    .S(_03235_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_1 _19191_ (.A(_03238_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_2 _19192_ (.A0(\core.cpuregs[14][5] ),
    .A1(_03101_),
    .S(_03235_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_1 _19193_ (.A(_03239_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _19194_ (.A0(\core.cpuregs[14][6] ),
    .A1(_03103_),
    .S(_03235_),
    .X(_03240_));
 sky130_fd_sc_hd__clkbuf_1 _19195_ (.A(_03240_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _19196_ (.A0(\core.cpuregs[14][7] ),
    .A1(_03105_),
    .S(_03235_),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_8 _19197_ (.A(_03241_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _19198_ (.A0(\core.cpuregs[14][8] ),
    .A1(_03107_),
    .S(_03231_),
    .X(_03242_));
 sky130_fd_sc_hd__clkbuf_1 _19199_ (.A(_03242_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _19200_ (.A0(\core.cpuregs[14][9] ),
    .A1(_03109_),
    .S(_03231_),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_1 _19201_ (.A(_03243_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19202_ (.A0(\core.cpuregs[14][10] ),
    .A1(_03111_),
    .S(_03231_),
    .X(_03244_));
 sky130_fd_sc_hd__clkbuf_1 _19203_ (.A(_03244_),
    .X(_00905_));
 sky130_fd_sc_hd__inv_2 _19204_ (.A(_03230_),
    .Y(_03245_));
 sky130_fd_sc_hd__clkbuf_2 _19205_ (.A(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _19206_ (.A0(_03113_),
    .A1(\core.cpuregs[14][11] ),
    .S(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__clkbuf_1 _19207_ (.A(_03247_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19208_ (.A0(\core.cpuregs[14][12] ),
    .A1(_03117_),
    .S(_03231_),
    .X(_03248_));
 sky130_fd_sc_hd__clkbuf_1 _19209_ (.A(_03248_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19210_ (.A0(_03119_),
    .A1(\core.cpuregs[14][13] ),
    .S(_03246_),
    .X(_03249_));
 sky130_fd_sc_hd__clkbuf_2 _19211_ (.A(_03249_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_8 _19212_ (.A0(_03121_),
    .A1(\core.cpuregs[14][14] ),
    .S(_03245_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_1 _19213_ (.A(_03250_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _19214_ (.A0(_03123_),
    .A1(\core.cpuregs[14][15] ),
    .S(_03245_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_1 _19215_ (.A(_03251_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _19216_ (.A0(_03125_),
    .A1(\core.cpuregs[14][16] ),
    .S(_03245_),
    .X(_03252_));
 sky130_fd_sc_hd__clkbuf_1 _19217_ (.A(_03252_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19218_ (.A0(_03127_),
    .A1(\core.cpuregs[14][17] ),
    .S(_03245_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_1 _19219_ (.A(_03253_),
    .X(_00912_));
 sky130_fd_sc_hd__nand2_1 _19220_ (.A(_03246_),
    .B(\core.cpuregs[14][18] ),
    .Y(_03254_));
 sky130_fd_sc_hd__a21bo_1 _19221_ (.A1(_03198_),
    .A2(_03232_),
    .B1_N(_03254_),
    .X(_00913_));
 sky130_fd_sc_hd__clkbuf_4 _19222_ (.A(_03232_),
    .X(_03255_));
 sky130_fd_sc_hd__nand2_1 _19223_ (.A(_03130_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__clkbuf_4 _19224_ (.A(_03246_),
    .X(_03257_));
 sky130_fd_sc_hd__nand2_1 _19225_ (.A(_03257_),
    .B(\core.cpuregs[14][19] ),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_1 _19226_ (.A(_03256_),
    .B(_03258_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _19227_ (.A(_03135_),
    .B(_03255_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _19228_ (.A(_03257_),
    .B(\core.cpuregs[14][20] ),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_1 _19229_ (.A(_03259_),
    .B(_03260_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_1 _19230_ (.A(_03138_),
    .B(_03255_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand2_1 _19231_ (.A(_03257_),
    .B(\core.cpuregs[14][21] ),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _19232_ (.A(_03261_),
    .B(_03262_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand2_1 _19233_ (.A(_03141_),
    .B(_03255_),
    .Y(_03263_));
 sky130_fd_sc_hd__nand2_1 _19234_ (.A(_03257_),
    .B(\core.cpuregs[14][22] ),
    .Y(_03264_));
 sky130_fd_sc_hd__nand2_1 _19235_ (.A(_03263_),
    .B(_03264_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _19236_ (.A(_03144_),
    .B(_03255_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _19237_ (.A(_03257_),
    .B(\core.cpuregs[14][23] ),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _19238_ (.A(_03265_),
    .B(_03266_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_1 _19239_ (.A(_03147_),
    .B(_03255_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_1 _19240_ (.A(_03257_),
    .B(\core.cpuregs[14][24] ),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _19241_ (.A(_03267_),
    .B(_03268_),
    .Y(_00919_));
 sky130_fd_sc_hd__clkbuf_2 _19242_ (.A(_03232_),
    .X(_03269_));
 sky130_fd_sc_hd__nand2_1 _19243_ (.A(_03150_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19244_ (.A(_03246_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2_1 _19245_ (.A(_03271_),
    .B(net131),
    .Y(_03272_));
 sky130_fd_sc_hd__nand2_1 _19246_ (.A(_03270_),
    .B(_03272_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_1 _19247_ (.A(_03155_),
    .B(_03269_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_1 _19248_ (.A(_03271_),
    .B(net142),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _19249_ (.A(_03273_),
    .B(_03274_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand2_1 _19250_ (.A(_03158_),
    .B(_03269_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _19251_ (.A(_03271_),
    .B(\core.cpuregs[14][27] ),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _19252_ (.A(_03275_),
    .B(_03276_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_1 _19253_ (.A(_03161_),
    .B(_03269_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_2 _19254_ (.A(_03271_),
    .B(\core.cpuregs[14][28] ),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _19255_ (.A(_03277_),
    .B(_03278_),
    .Y(_00923_));
 sky130_fd_sc_hd__nand2_4 _19256_ (.A(_03164_),
    .B(_03269_),
    .Y(_03279_));
 sky130_fd_sc_hd__nand2_1 _19257_ (.A(_03271_),
    .B(\core.cpuregs[14][29] ),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _19258_ (.A(_03279_),
    .B(_03280_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _19259_ (.A(_03167_),
    .B(_03269_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _19260_ (.A(_03271_),
    .B(\core.cpuregs[14][30] ),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _19261_ (.A(_03281_),
    .B(_03282_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _19262_ (.A(_03170_),
    .B(_03232_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand2_1 _19263_ (.A(_03246_),
    .B(net139),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _19264_ (.A(_03283_),
    .B(_03284_),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _19265_ (.A(_03173_),
    .B(_02778_),
    .Y(_03285_));
 sky130_fd_sc_hd__clkbuf_4 _19266_ (.A(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__clkbuf_2 _19267_ (.A(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__mux2_2 _19268_ (.A0(\core.cpuregs[13][0] ),
    .A1(_03087_),
    .S(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_1 _19269_ (.A(_03288_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19270_ (.A0(\core.cpuregs[13][1] ),
    .A1(_03092_),
    .S(_03287_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_1 _19271_ (.A(_03289_),
    .X(_00928_));
 sky130_fd_sc_hd__clkbuf_4 _19272_ (.A(_03286_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _19273_ (.A0(\core.cpuregs[13][2] ),
    .A1(_03094_),
    .S(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_4 _19274_ (.A(_03291_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19275_ (.A0(\core.cpuregs[13][3] ),
    .A1(_03097_),
    .S(_03290_),
    .X(_03292_));
 sky130_fd_sc_hd__buf_1 _19276_ (.A(_03292_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19277_ (.A0(\core.cpuregs[13][4] ),
    .A1(_03099_),
    .S(_03290_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_1 _19278_ (.A(_03293_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_2 _19279_ (.A0(\core.cpuregs[13][5] ),
    .A1(_03101_),
    .S(_03290_),
    .X(_03294_));
 sky130_fd_sc_hd__clkbuf_1 _19280_ (.A(_03294_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19281_ (.A0(\core.cpuregs[13][6] ),
    .A1(_03103_),
    .S(_03290_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_1 _19282_ (.A(_03295_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19283_ (.A0(\core.cpuregs[13][7] ),
    .A1(_03105_),
    .S(_03290_),
    .X(_03296_));
 sky130_fd_sc_hd__clkbuf_1 _19284_ (.A(_03296_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _19285_ (.A0(\core.cpuregs[13][8] ),
    .A1(_03107_),
    .S(_03286_),
    .X(_03297_));
 sky130_fd_sc_hd__clkbuf_1 _19286_ (.A(_03297_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _19287_ (.A0(\core.cpuregs[13][9] ),
    .A1(_03109_),
    .S(_03286_),
    .X(_03298_));
 sky130_fd_sc_hd__clkbuf_2 _19288_ (.A(_03298_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19289_ (.A0(\core.cpuregs[13][10] ),
    .A1(_03111_),
    .S(_03286_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_1 _19290_ (.A(_03299_),
    .X(_00937_));
 sky130_fd_sc_hd__inv_2 _19291_ (.A(_03285_),
    .Y(_03300_));
 sky130_fd_sc_hd__clkbuf_4 _19292_ (.A(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _19293_ (.A0(_03113_),
    .A1(\core.cpuregs[13][11] ),
    .S(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_1 _19294_ (.A(_03302_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19295_ (.A0(\core.cpuregs[13][12] ),
    .A1(_03117_),
    .S(_03286_),
    .X(_03303_));
 sky130_fd_sc_hd__clkbuf_1 _19296_ (.A(_03303_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19297_ (.A0(_03119_),
    .A1(\core.cpuregs[13][13] ),
    .S(_03301_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_1 _19298_ (.A(_03304_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19299_ (.A0(_03121_),
    .A1(\core.cpuregs[13][14] ),
    .S(_03300_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_2 _19300_ (.A(_03305_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _19301_ (.A0(_03123_),
    .A1(\core.cpuregs[13][15] ),
    .S(_03300_),
    .X(_03306_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19302_ (.A(_03306_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_4 _19303_ (.A0(_03125_),
    .A1(\core.cpuregs[13][16] ),
    .S(_03300_),
    .X(_03307_));
 sky130_fd_sc_hd__clkbuf_1 _19304_ (.A(_03307_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _19305_ (.A0(_03127_),
    .A1(\core.cpuregs[13][17] ),
    .S(_03300_),
    .X(_03308_));
 sky130_fd_sc_hd__clkbuf_2 _19306_ (.A(_03308_),
    .X(_00944_));
 sky130_fd_sc_hd__nand2_1 _19307_ (.A(_03301_),
    .B(\core.cpuregs[13][18] ),
    .Y(_03309_));
 sky130_fd_sc_hd__a21bo_1 _19308_ (.A1(_03198_),
    .A2(_03287_),
    .B1_N(_03309_),
    .X(_00945_));
 sky130_fd_sc_hd__clkbuf_4 _19309_ (.A(_03287_),
    .X(_03310_));
 sky130_fd_sc_hd__nand2_1 _19310_ (.A(_03130_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__buf_2 _19311_ (.A(_03301_),
    .X(_03312_));
 sky130_fd_sc_hd__nand2_1 _19312_ (.A(_03312_),
    .B(\core.cpuregs[13][19] ),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(_03311_),
    .B(_03313_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _19314_ (.A(_03135_),
    .B(_03310_),
    .Y(_03314_));
 sky130_fd_sc_hd__nand2_1 _19315_ (.A(_03312_),
    .B(\core.cpuregs[13][20] ),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _19316_ (.A(_03314_),
    .B(_03315_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _19317_ (.A(_03138_),
    .B(_03310_),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _19318_ (.A(_03312_),
    .B(net160),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_1 _19319_ (.A(_03316_),
    .B(_03317_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _19320_ (.A(_03141_),
    .B(_03310_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _19321_ (.A(_03312_),
    .B(net167),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2_1 _19322_ (.A(_03318_),
    .B(_03319_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _19323_ (.A(_03144_),
    .B(_03310_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _19324_ (.A(_03312_),
    .B(\core.cpuregs[13][23] ),
    .Y(_03321_));
 sky130_fd_sc_hd__nand2_1 _19325_ (.A(_03320_),
    .B(_03321_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2_1 _19326_ (.A(_03147_),
    .B(_03310_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _19327_ (.A(_03312_),
    .B(net132),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _19328_ (.A(_03322_),
    .B(_03323_),
    .Y(_00951_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19329_ (.A(_03287_),
    .X(_03324_));
 sky130_fd_sc_hd__nand2_1 _19330_ (.A(_03150_),
    .B(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19331_ (.A(_03301_),
    .X(_03326_));
 sky130_fd_sc_hd__nand2_1 _19332_ (.A(_03326_),
    .B(\core.cpuregs[13][25] ),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_03325_),
    .B(_03327_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _19334_ (.A(_03155_),
    .B(_03324_),
    .Y(_03328_));
 sky130_fd_sc_hd__nand2_1 _19335_ (.A(_03326_),
    .B(\core.cpuregs[13][26] ),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _19336_ (.A(_03328_),
    .B(_03329_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _19337_ (.A(_03158_),
    .B(_03324_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _19338_ (.A(_03326_),
    .B(\core.cpuregs[13][27] ),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _19339_ (.A(_03330_),
    .B(_03331_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand2_1 _19340_ (.A(_03161_),
    .B(_03324_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_1 _19341_ (.A(_03326_),
    .B(\core.cpuregs[13][28] ),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _19342_ (.A(_03332_),
    .B(_03333_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _19343_ (.A(_03164_),
    .B(_03324_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand2_1 _19344_ (.A(_03326_),
    .B(\core.cpuregs[13][29] ),
    .Y(_03335_));
 sky130_fd_sc_hd__nand2_1 _19345_ (.A(_03334_),
    .B(_03335_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2_1 _19346_ (.A(_03167_),
    .B(_03324_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _19347_ (.A(_03326_),
    .B(\core.cpuregs[13][30] ),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _19348_ (.A(_03336_),
    .B(_03337_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_2 _19349_ (.A(_03170_),
    .B(_03287_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_2 _19350_ (.A(_03301_),
    .B(\core.cpuregs[13][31] ),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_8 _19351_ (.A(_03338_),
    .B(_03339_),
    .Y(_00958_));
 sky130_fd_sc_hd__nor2_8 _19352_ (.A(_03173_),
    .B(_09950_),
    .Y(_03340_));
 sky130_fd_sc_hd__clkbuf_4 _19353_ (.A(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_2 _19354_ (.A(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_2 _19355_ (.A0(\core.cpuregs[12][0] ),
    .A1(_03087_),
    .S(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _19356_ (.A(_03343_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19357_ (.A0(\core.cpuregs[12][1] ),
    .A1(_03092_),
    .S(_03342_),
    .X(_03344_));
 sky130_fd_sc_hd__clkbuf_1 _19358_ (.A(_03344_),
    .X(_00960_));
 sky130_fd_sc_hd__clkbuf_4 _19359_ (.A(_03341_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _19360_ (.A0(\core.cpuregs[12][2] ),
    .A1(_03094_),
    .S(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__buf_1 _19361_ (.A(_03346_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _19362_ (.A0(\core.cpuregs[12][3] ),
    .A1(_03097_),
    .S(_03345_),
    .X(_03347_));
 sky130_fd_sc_hd__buf_1 _19363_ (.A(_03347_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _19364_ (.A0(\core.cpuregs[12][4] ),
    .A1(_03099_),
    .S(_03345_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _19365_ (.A(_03348_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_2 _19366_ (.A0(\core.cpuregs[12][5] ),
    .A1(_03101_),
    .S(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__clkbuf_4 _19367_ (.A(_03349_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _19368_ (.A0(\core.cpuregs[12][6] ),
    .A1(_03103_),
    .S(_03345_),
    .X(_03350_));
 sky130_fd_sc_hd__clkbuf_1 _19369_ (.A(_03350_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _19370_ (.A0(\core.cpuregs[12][7] ),
    .A1(_03105_),
    .S(_03345_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_4 _19371_ (.A(_03351_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19372_ (.A0(\core.cpuregs[12][8] ),
    .A1(_03107_),
    .S(_03341_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_4 _19373_ (.A(_03352_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19374_ (.A0(\core.cpuregs[12][9] ),
    .A1(_03109_),
    .S(_03341_),
    .X(_03353_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19375_ (.A(_03353_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _19376_ (.A0(\core.cpuregs[12][10] ),
    .A1(_03111_),
    .S(_03341_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _19377_ (.A(_03354_),
    .X(_00969_));
 sky130_fd_sc_hd__inv_2 _19378_ (.A(_03340_),
    .Y(_03355_));
 sky130_fd_sc_hd__clkbuf_4 _19379_ (.A(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _19380_ (.A0(_03113_),
    .A1(\core.cpuregs[12][11] ),
    .S(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _19381_ (.A(_03357_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _19382_ (.A0(\core.cpuregs[12][12] ),
    .A1(_03117_),
    .S(_03341_),
    .X(_03358_));
 sky130_fd_sc_hd__clkbuf_8 _19383_ (.A(_03358_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19384_ (.A0(_03119_),
    .A1(\core.cpuregs[12][13] ),
    .S(_03356_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _19385_ (.A(_03359_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19386_ (.A0(_03121_),
    .A1(\core.cpuregs[12][14] ),
    .S(_03355_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_2 _19387_ (.A(_03360_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _19388_ (.A0(_03123_),
    .A1(\core.cpuregs[12][15] ),
    .S(_03355_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_1 _19389_ (.A(_03361_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_4 _19390_ (.A0(_03125_),
    .A1(\core.cpuregs[12][16] ),
    .S(_03355_),
    .X(_03362_));
 sky130_fd_sc_hd__clkbuf_1 _19391_ (.A(_03362_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _19392_ (.A0(_03127_),
    .A1(\core.cpuregs[12][17] ),
    .S(_03355_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_2 _19393_ (.A(_03363_),
    .X(_00976_));
 sky130_fd_sc_hd__nand2_1 _19394_ (.A(_03356_),
    .B(\core.cpuregs[12][18] ),
    .Y(_03364_));
 sky130_fd_sc_hd__a21bo_1 _19395_ (.A1(_03198_),
    .A2(_03342_),
    .B1_N(_03364_),
    .X(_00977_));
 sky130_fd_sc_hd__clkbuf_4 _19396_ (.A(_03342_),
    .X(_03365_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(_03130_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__buf_2 _19398_ (.A(_03356_),
    .X(_03367_));
 sky130_fd_sc_hd__nand2_1 _19399_ (.A(_03367_),
    .B(net141),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _19400_ (.A(_03366_),
    .B(_03368_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_1 _19401_ (.A(_03135_),
    .B(_03365_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _19402_ (.A(_03367_),
    .B(\core.cpuregs[12][20] ),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_1 _19403_ (.A(_03369_),
    .B(_03370_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _19404_ (.A(_03138_),
    .B(_03365_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _19405_ (.A(_03367_),
    .B(\core.cpuregs[12][21] ),
    .Y(_03372_));
 sky130_fd_sc_hd__nand2_1 _19406_ (.A(_03371_),
    .B(_03372_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _19407_ (.A(_03141_),
    .B(_03365_),
    .Y(_03373_));
 sky130_fd_sc_hd__nand2_1 _19408_ (.A(_03367_),
    .B(\core.cpuregs[12][22] ),
    .Y(_03374_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(_03373_),
    .B(_03374_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _19410_ (.A(_03144_),
    .B(_03365_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand2_1 _19411_ (.A(_03367_),
    .B(\core.cpuregs[12][23] ),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _19412_ (.A(_03375_),
    .B(_03376_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _19413_ (.A(_03147_),
    .B(_03365_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _19414_ (.A(_03367_),
    .B(net144),
    .Y(_03378_));
 sky130_fd_sc_hd__nand2_1 _19415_ (.A(_03377_),
    .B(_03378_),
    .Y(_00983_));
 sky130_fd_sc_hd__clkbuf_2 _19416_ (.A(_03342_),
    .X(_03379_));
 sky130_fd_sc_hd__nand2_1 _19417_ (.A(_03150_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__clkbuf_4 _19418_ (.A(_03356_),
    .X(_03381_));
 sky130_fd_sc_hd__nand2_1 _19419_ (.A(_03381_),
    .B(\core.cpuregs[12][25] ),
    .Y(_03382_));
 sky130_fd_sc_hd__nand2_1 _19420_ (.A(_03380_),
    .B(_03382_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _19421_ (.A(_03155_),
    .B(_03379_),
    .Y(_03383_));
 sky130_fd_sc_hd__nand2_1 _19422_ (.A(_03381_),
    .B(net137),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _19423_ (.A(_03383_),
    .B(_03384_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _19424_ (.A(_03158_),
    .B(_03379_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2_1 _19425_ (.A(_03381_),
    .B(\core.cpuregs[12][27] ),
    .Y(_03386_));
 sky130_fd_sc_hd__nand2_1 _19426_ (.A(_03385_),
    .B(_03386_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _19427_ (.A(_03161_),
    .B(_03379_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _19428_ (.A(_03381_),
    .B(net130),
    .Y(_03388_));
 sky130_fd_sc_hd__nand2_1 _19429_ (.A(_03387_),
    .B(_03388_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _19430_ (.A(_03164_),
    .B(_03379_),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _19431_ (.A(_03381_),
    .B(net170),
    .Y(_03390_));
 sky130_fd_sc_hd__nand2_1 _19432_ (.A(_03389_),
    .B(_03390_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _19433_ (.A(_03167_),
    .B(_03379_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _19434_ (.A(_03381_),
    .B(\core.cpuregs[12][30] ),
    .Y(_03392_));
 sky130_fd_sc_hd__nand2_1 _19435_ (.A(_03391_),
    .B(_03392_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _19436_ (.A(_03170_),
    .B(_03342_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _19437_ (.A(_03356_),
    .B(\core.cpuregs[12][31] ),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _19438_ (.A(_03393_),
    .B(_03394_),
    .Y(_00990_));
 sky130_fd_sc_hd__and3_1 _19439_ (.A(_09317_),
    .B(_09319_),
    .C(\core.latched_rd[3] ),
    .X(_03395_));
 sky130_fd_sc_hd__inv_2 _19440_ (.A(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nor2_1 _19441_ (.A(_03396_),
    .B(_09812_),
    .Y(_03397_));
 sky130_fd_sc_hd__clkbuf_4 _19442_ (.A(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _19443_ (.A0(\core.cpuregs[11][0] ),
    .A1(_03087_),
    .S(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _19444_ (.A(_03399_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _19445_ (.A0(\core.cpuregs[11][1] ),
    .A1(_03092_),
    .S(_03398_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _19446_ (.A(_03400_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _19447_ (.A0(\core.cpuregs[11][2] ),
    .A1(_03094_),
    .S(_03398_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _19448_ (.A(_03401_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _19449_ (.A0(\core.cpuregs[11][3] ),
    .A1(_03097_),
    .S(_03398_),
    .X(_03402_));
 sky130_fd_sc_hd__buf_1 _19450_ (.A(_03402_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _19451_ (.A0(\core.cpuregs[11][4] ),
    .A1(_03099_),
    .S(_03398_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _19452_ (.A(_03403_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_2 _19453_ (.A0(\core.cpuregs[11][5] ),
    .A1(_03101_),
    .S(_03398_),
    .X(_03404_));
 sky130_fd_sc_hd__buf_4 _19454_ (.A(_03404_),
    .X(_00996_));
 sky130_fd_sc_hd__clkbuf_2 _19455_ (.A(_03397_),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_2 _19456_ (.A0(\core.cpuregs[11][6] ),
    .A1(_03103_),
    .S(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__buf_4 _19457_ (.A(_03406_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _19458_ (.A0(\core.cpuregs[11][7] ),
    .A1(_03105_),
    .S(_03405_),
    .X(_03407_));
 sky130_fd_sc_hd__buf_4 _19459_ (.A(_03407_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_4 _19460_ (.A0(\core.cpuregs[11][8] ),
    .A1(_03107_),
    .S(_03405_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(_03408_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_2 _19462_ (.A0(\core.cpuregs[11][9] ),
    .A1(_03109_),
    .S(_03405_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _19463_ (.A(_03409_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _19464_ (.A0(\core.cpuregs[11][10] ),
    .A1(_03111_),
    .S(_03405_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _19465_ (.A(_03410_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _19466_ (.A(_09324_),
    .B(_09326_),
    .C(_03395_),
    .X(_03411_));
 sky130_fd_sc_hd__inv_2 _19467_ (.A(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__clkbuf_2 _19468_ (.A(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_8 _19469_ (.A0(_03113_),
    .A1(\core.cpuregs[11][11] ),
    .S(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _19470_ (.A(_03414_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _19471_ (.A0(\core.cpuregs[11][12] ),
    .A1(_03117_),
    .S(_03405_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_4 _19472_ (.A(_03415_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _19473_ (.A0(_03119_),
    .A1(\core.cpuregs[11][13] ),
    .S(_03413_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _19474_ (.A(_03416_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _19475_ (.A0(_03121_),
    .A1(\core.cpuregs[11][14] ),
    .S(_03413_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _19476_ (.A(_03417_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _19477_ (.A0(_03123_),
    .A1(\core.cpuregs[11][15] ),
    .S(_03413_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _19478_ (.A(_03418_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_2 _19479_ (.A0(_03125_),
    .A1(\core.cpuregs[11][16] ),
    .S(_03413_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _19480_ (.A(_03419_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _19481_ (.A0(_03127_),
    .A1(\core.cpuregs[11][17] ),
    .S(_03412_),
    .X(_03420_));
 sky130_fd_sc_hd__clkbuf_8 _19482_ (.A(_03420_),
    .X(_01008_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19483_ (.A(_03397_),
    .X(_03421_));
 sky130_fd_sc_hd__and2_1 _19484_ (.A(_03413_),
    .B(\core.cpuregs[11][18] ),
    .X(_03422_));
 sky130_fd_sc_hd__a21o_1 _19485_ (.A1(_09779_),
    .A2(_03421_),
    .B1(_03422_),
    .X(_01009_));
 sky130_fd_sc_hd__inv_2 _19486_ (.A(\core.cpuregs[11][19] ),
    .Y(_03423_));
 sky130_fd_sc_hd__buf_4 _19487_ (.A(_09447_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_2 _19488_ (.A(_03421_),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_1 _19489_ (.A(_03424_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__o21ai_1 _19490_ (.A1(_03423_),
    .A2(_03421_),
    .B1(_03426_),
    .Y(_01010_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19491_ (.A(_03421_),
    .X(_03427_));
 sky130_fd_sc_hd__nand2_1 _19492_ (.A(_03135_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19493_ (.A(_03412_),
    .X(_03429_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19494_ (.A(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_1 _19495_ (.A(_03430_),
    .B(\core.cpuregs[11][20] ),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _19496_ (.A(_03428_),
    .B(_03431_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _19497_ (.A(_03138_),
    .B(_03427_),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2_1 _19498_ (.A(_03430_),
    .B(\core.cpuregs[11][21] ),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _19499_ (.A(_03432_),
    .B(_03433_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _19500_ (.A(\core.cpuregs[11][22] ),
    .Y(_03434_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19501_ (.A(_09473_),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_1 _19502_ (.A(_03435_),
    .B(_03421_),
    .Y(_03436_));
 sky130_fd_sc_hd__o21ai_1 _19503_ (.A1(_03434_),
    .A2(_03421_),
    .B1(_03436_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _19504_ (.A(_03144_),
    .B(_03427_),
    .Y(_03437_));
 sky130_fd_sc_hd__nand2_1 _19505_ (.A(_03430_),
    .B(\core.cpuregs[11][23] ),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_1 _19506_ (.A(_03437_),
    .B(_03438_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _19507_ (.A(_03147_),
    .B(_03427_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2_1 _19508_ (.A(_03430_),
    .B(\core.cpuregs[11][24] ),
    .Y(_03440_));
 sky130_fd_sc_hd__nand2_1 _19509_ (.A(_03439_),
    .B(_03440_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _19510_ (.A(_03150_),
    .B(_03427_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _19511_ (.A(_03430_),
    .B(\core.cpuregs[11][25] ),
    .Y(_03442_));
 sky130_fd_sc_hd__nand2_1 _19512_ (.A(_03441_),
    .B(_03442_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _19513_ (.A(_03155_),
    .B(_03427_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_1 _19514_ (.A(_03430_),
    .B(\core.cpuregs[11][26] ),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _19515_ (.A(_03443_),
    .B(_03444_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _19516_ (.A(_03158_),
    .B(_03425_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand2_1 _19517_ (.A(_03429_),
    .B(net183),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _19518_ (.A(_03445_),
    .B(_03446_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _19519_ (.A(_03161_),
    .B(_03425_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _19520_ (.A(_03429_),
    .B(\core.cpuregs[11][28] ),
    .Y(_03448_));
 sky130_fd_sc_hd__nand2_1 _19521_ (.A(_03447_),
    .B(_03448_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_2 _19522_ (.A(_03164_),
    .B(_03425_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _19523_ (.A(_03429_),
    .B(\core.cpuregs[11][29] ),
    .Y(_03450_));
 sky130_fd_sc_hd__nand2_1 _19524_ (.A(_03449_),
    .B(_03450_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_2 _19525_ (.A(_03167_),
    .B(_03425_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_1 _19526_ (.A(_03429_),
    .B(\core.cpuregs[11][30] ),
    .Y(_03452_));
 sky130_fd_sc_hd__nand2_1 _19527_ (.A(_03451_),
    .B(_03452_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _19528_ (.A(_03170_),
    .B(_03425_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand2_1 _19529_ (.A(_03429_),
    .B(\core.cpuregs[11][31] ),
    .Y(_03454_));
 sky130_fd_sc_hd__nand2_1 _19530_ (.A(_03453_),
    .B(_03454_),
    .Y(_01022_));
 sky130_fd_sc_hd__buf_1 _19531_ (.A(_09314_),
    .X(_03455_));
 sky130_fd_sc_hd__nor2_1 _19532_ (.A(_03396_),
    .B(_10158_),
    .Y(_03456_));
 sky130_fd_sc_hd__clkbuf_4 _19533_ (.A(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__mux2_1 _19534_ (.A0(\core.cpuregs[10][0] ),
    .A1(_03455_),
    .S(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_1 _19535_ (.A(_03458_),
    .X(_01023_));
 sky130_fd_sc_hd__buf_1 _19536_ (.A(_09336_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2_1 _19537_ (.A0(\core.cpuregs[10][1] ),
    .A1(_03459_),
    .S(_03457_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_1 _19538_ (.A(_03460_),
    .X(_01024_));
 sky130_fd_sc_hd__buf_2 _19539_ (.A(_09339_),
    .X(_03461_));
 sky130_fd_sc_hd__mux2_1 _19540_ (.A0(\core.cpuregs[10][2] ),
    .A1(_03461_),
    .S(_03457_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_1 _19541_ (.A(_03462_),
    .X(_01025_));
 sky130_fd_sc_hd__buf_2 _19542_ (.A(_09348_),
    .X(_03463_));
 sky130_fd_sc_hd__mux2_1 _19543_ (.A0(\core.cpuregs[10][3] ),
    .A1(_03463_),
    .S(_03457_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_2 _19544_ (.A(_03464_),
    .X(_01026_));
 sky130_fd_sc_hd__buf_2 _19545_ (.A(_09356_),
    .X(_03465_));
 sky130_fd_sc_hd__mux2_1 _19546_ (.A0(\core.cpuregs[10][4] ),
    .A1(_03465_),
    .S(_03457_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_1 _19547_ (.A(_03466_),
    .X(_01027_));
 sky130_fd_sc_hd__clkbuf_2 _19548_ (.A(_09362_),
    .X(_03467_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(\core.cpuregs[10][5] ),
    .A1(_03467_),
    .S(_03457_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _19550_ (.A(_03468_),
    .X(_01028_));
 sky130_fd_sc_hd__buf_2 _19551_ (.A(_09368_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_2 _19552_ (.A(_03456_),
    .X(_03470_));
 sky130_fd_sc_hd__mux2_1 _19553_ (.A0(\core.cpuregs[10][6] ),
    .A1(_03469_),
    .S(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _19554_ (.A(_03471_),
    .X(_01029_));
 sky130_fd_sc_hd__buf_1 _19555_ (.A(_09374_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _19556_ (.A0(\core.cpuregs[10][7] ),
    .A1(_03472_),
    .S(_03470_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _19557_ (.A(_03473_),
    .X(_01030_));
 sky130_fd_sc_hd__buf_1 _19558_ (.A(_09380_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _19559_ (.A0(\core.cpuregs[10][8] ),
    .A1(_03474_),
    .S(_03470_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _19560_ (.A(_03475_),
    .X(_01031_));
 sky130_fd_sc_hd__buf_1 _19561_ (.A(_09387_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_2 _19562_ (.A0(\core.cpuregs[10][9] ),
    .A1(_03476_),
    .S(_03470_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _19563_ (.A(_03477_),
    .X(_01032_));
 sky130_fd_sc_hd__clkbuf_4 _19564_ (.A(_09394_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _19565_ (.A0(\core.cpuregs[10][10] ),
    .A1(_03478_),
    .S(_03470_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_1 _19566_ (.A(_03479_),
    .X(_01033_));
 sky130_fd_sc_hd__buf_1 _19567_ (.A(_09400_),
    .X(_03480_));
 sky130_fd_sc_hd__and3_4 _19568_ (.A(_09324_),
    .B(_09556_),
    .C(_03395_),
    .X(_03481_));
 sky130_fd_sc_hd__inv_2 _19569_ (.A(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__clkbuf_2 _19570_ (.A(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_8 _19571_ (.A0(_03480_),
    .A1(\core.cpuregs[10][11] ),
    .S(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _19572_ (.A(_03484_),
    .X(_01034_));
 sky130_fd_sc_hd__clkbuf_4 _19573_ (.A(_09407_),
    .X(_03485_));
 sky130_fd_sc_hd__mux2_1 _19574_ (.A0(\core.cpuregs[10][12] ),
    .A1(_03485_),
    .S(_03470_),
    .X(_03486_));
 sky130_fd_sc_hd__buf_4 _19575_ (.A(_03486_),
    .X(_01035_));
 sky130_fd_sc_hd__buf_2 _19576_ (.A(_09413_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _19577_ (.A0(_03487_),
    .A1(\core.cpuregs[10][13] ),
    .S(_03483_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _19578_ (.A(_03488_),
    .X(_01036_));
 sky130_fd_sc_hd__buf_1 _19579_ (.A(_09418_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _19580_ (.A0(_03489_),
    .A1(\core.cpuregs[10][14] ),
    .S(_03483_),
    .X(_03490_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19581_ (.A(_03490_),
    .X(_01037_));
 sky130_fd_sc_hd__clkbuf_2 _19582_ (.A(_09423_),
    .X(_03491_));
 sky130_fd_sc_hd__mux2_1 _19583_ (.A0(_03491_),
    .A1(\core.cpuregs[10][15] ),
    .S(_03483_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _19584_ (.A(_03492_),
    .X(_01038_));
 sky130_fd_sc_hd__buf_1 _19585_ (.A(_09430_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_4 _19586_ (.A0(_03493_),
    .A1(\core.cpuregs[10][16] ),
    .S(_03483_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _19587_ (.A(_03494_),
    .X(_01039_));
 sky130_fd_sc_hd__buf_2 _19588_ (.A(_09435_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _19589_ (.A0(_03495_),
    .A1(\core.cpuregs[10][17] ),
    .S(_03482_),
    .X(_03496_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19590_ (.A(_03496_),
    .X(_01040_));
 sky130_fd_sc_hd__clkbuf_2 _19591_ (.A(_03456_),
    .X(_03497_));
 sky130_fd_sc_hd__and2_1 _19592_ (.A(_03483_),
    .B(\core.cpuregs[10][18] ),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _19593_ (.A1(_09779_),
    .A2(_03497_),
    .B1(_03498_),
    .X(_01041_));
 sky130_fd_sc_hd__inv_2 _19594_ (.A(\core.cpuregs[10][19] ),
    .Y(_03499_));
 sky130_fd_sc_hd__buf_2 _19595_ (.A(_03497_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_1 _19596_ (.A(_03424_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__o21ai_2 _19597_ (.A1(_03499_),
    .A2(_03497_),
    .B1(_03501_),
    .Y(_01042_));
 sky130_fd_sc_hd__clkbuf_2 _19598_ (.A(_09457_),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_2 _19599_ (.A(_03497_),
    .X(_03503_));
 sky130_fd_sc_hd__nand2_2 _19600_ (.A(_03502_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__clkbuf_4 _19601_ (.A(_03482_),
    .X(_03505_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19602_ (.A(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__nand2_1 _19603_ (.A(_03506_),
    .B(\core.cpuregs[10][20] ),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(_03504_),
    .B(_03507_),
    .Y(_01043_));
 sky130_fd_sc_hd__buf_6 _19605_ (.A(_09466_),
    .X(_03508_));
 sky130_fd_sc_hd__nand2_4 _19606_ (.A(_03508_),
    .B(_03503_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand2_1 _19607_ (.A(_03506_),
    .B(\core.cpuregs[10][21] ),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_4 _19608_ (.A(_03509_),
    .B(_03510_),
    .Y(_01044_));
 sky130_fd_sc_hd__inv_2 _19609_ (.A(net174),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _19610_ (.A(_03435_),
    .B(_03497_),
    .Y(_03512_));
 sky130_fd_sc_hd__o21ai_1 _19611_ (.A1(_03511_),
    .A2(_03497_),
    .B1(_03512_),
    .Y(_01045_));
 sky130_fd_sc_hd__buf_6 _19612_ (.A(_09480_),
    .X(_03513_));
 sky130_fd_sc_hd__nand2_1 _19613_ (.A(_03513_),
    .B(_03503_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_03506_),
    .B(net156),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _19615_ (.A(_03514_),
    .B(_03515_),
    .Y(_01046_));
 sky130_fd_sc_hd__buf_6 _19616_ (.A(_09488_),
    .X(_03516_));
 sky130_fd_sc_hd__nand2_1 _19617_ (.A(_03516_),
    .B(_03503_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _19618_ (.A(_03506_),
    .B(net148),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_1 _19619_ (.A(_03517_),
    .B(_03518_),
    .Y(_01047_));
 sky130_fd_sc_hd__clkbuf_4 _19620_ (.A(_09498_),
    .X(_03519_));
 sky130_fd_sc_hd__nand2_1 _19621_ (.A(_03519_),
    .B(_03503_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _19622_ (.A(_03506_),
    .B(\core.cpuregs[10][25] ),
    .Y(_03521_));
 sky130_fd_sc_hd__nand2_1 _19623_ (.A(_03520_),
    .B(_03521_),
    .Y(_01048_));
 sky130_fd_sc_hd__clkbuf_2 _19624_ (.A(_09508_),
    .X(_03522_));
 sky130_fd_sc_hd__nand2_1 _19625_ (.A(_03522_),
    .B(_03503_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _19626_ (.A(_03506_),
    .B(\core.cpuregs[10][26] ),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_1 _19627_ (.A(_03523_),
    .B(_03524_),
    .Y(_01049_));
 sky130_fd_sc_hd__buf_6 _19628_ (.A(_09515_),
    .X(_03525_));
 sky130_fd_sc_hd__nand2_1 _19629_ (.A(_03525_),
    .B(_03500_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _19630_ (.A(_03505_),
    .B(net173),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _19631_ (.A(_03526_),
    .B(_03527_),
    .Y(_01050_));
 sky130_fd_sc_hd__buf_6 _19632_ (.A(_09524_),
    .X(_03528_));
 sky130_fd_sc_hd__nand2_1 _19633_ (.A(_03528_),
    .B(_03500_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _19634_ (.A(_03505_),
    .B(net123),
    .Y(_03530_));
 sky130_fd_sc_hd__nand2_1 _19635_ (.A(_03529_),
    .B(_03530_),
    .Y(_01051_));
 sky130_fd_sc_hd__buf_2 _19636_ (.A(_09533_),
    .X(_03531_));
 sky130_fd_sc_hd__nand2_1 _19637_ (.A(_03531_),
    .B(_03500_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2_1 _19638_ (.A(_03505_),
    .B(\core.cpuregs[10][29] ),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _19639_ (.A(_03532_),
    .B(_03533_),
    .Y(_01052_));
 sky130_fd_sc_hd__buf_6 _19640_ (.A(_09541_),
    .X(_03534_));
 sky130_fd_sc_hd__nand2_1 _19641_ (.A(_03534_),
    .B(_03500_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _19642_ (.A(_03505_),
    .B(\core.cpuregs[10][30] ),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _19643_ (.A(_03535_),
    .B(_03536_),
    .Y(_01053_));
 sky130_fd_sc_hd__buf_2 _19644_ (.A(_09550_),
    .X(_03537_));
 sky130_fd_sc_hd__nand2_1 _19645_ (.A(_03537_),
    .B(_03500_),
    .Y(_03538_));
 sky130_fd_sc_hd__nand2_1 _19646_ (.A(_03505_),
    .B(net140),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _19647_ (.A(_03538_),
    .B(_03539_),
    .Y(_01054_));
 sky130_fd_sc_hd__clkbuf_1 _19648_ (.A(\core.cpuregs[0][0] ),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_2 _19649_ (.A(_03540_),
    .X(_01055_));
 sky130_fd_sc_hd__clkbuf_1 _19650_ (.A(\core.cpuregs[0][1] ),
    .X(_03541_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19651_ (.A(_03541_),
    .X(_01056_));
 sky130_fd_sc_hd__buf_1 _19652_ (.A(\core.cpuregs[0][2] ),
    .X(_03542_));
 sky130_fd_sc_hd__buf_1 _19653_ (.A(_03542_),
    .X(_01057_));
 sky130_fd_sc_hd__buf_1 _19654_ (.A(\core.cpuregs[0][3] ),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _19655_ (.A(_03543_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_1 _19656_ (.A(\core.cpuregs[0][4] ),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _19657_ (.A(_03544_),
    .X(_01059_));
 sky130_fd_sc_hd__buf_2 _19658_ (.A(\core.cpuregs[0][5] ),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _19659_ (.A(_03545_),
    .X(_01060_));
 sky130_fd_sc_hd__buf_1 _19660_ (.A(\core.cpuregs[0][6] ),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _19661_ (.A(_03546_),
    .X(_01061_));
 sky130_fd_sc_hd__buf_1 _19662_ (.A(\core.cpuregs[0][7] ),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _19663_ (.A(_03547_),
    .X(_01062_));
 sky130_fd_sc_hd__buf_1 _19664_ (.A(\core.cpuregs[0][8] ),
    .X(_03548_));
 sky130_fd_sc_hd__buf_1 _19665_ (.A(_03548_),
    .X(_01063_));
 sky130_fd_sc_hd__clkbuf_1 _19666_ (.A(\core.cpuregs[0][9] ),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _19667_ (.A(_03549_),
    .X(_01064_));
 sky130_fd_sc_hd__clkbuf_2 _19668_ (.A(\core.cpuregs[0][10] ),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _19669_ (.A(_03550_),
    .X(_01065_));
 sky130_fd_sc_hd__clkbuf_1 _19670_ (.A(\core.cpuregs[0][11] ),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _19671_ (.A(_03551_),
    .X(_01066_));
 sky130_fd_sc_hd__clkbuf_1 _19672_ (.A(\core.cpuregs[0][12] ),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _19673_ (.A(_03552_),
    .X(_01067_));
 sky130_fd_sc_hd__buf_1 _19674_ (.A(\core.cpuregs[0][13] ),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _19675_ (.A(_03553_),
    .X(_01068_));
 sky130_fd_sc_hd__clkbuf_1 _19676_ (.A(\core.cpuregs[0][14] ),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _19677_ (.A(_03554_),
    .X(_01069_));
 sky130_fd_sc_hd__buf_1 _19678_ (.A(\core.cpuregs[0][15] ),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_2 _19679_ (.A(_03555_),
    .X(_01070_));
 sky130_fd_sc_hd__buf_1 _19680_ (.A(\core.cpuregs[0][16] ),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _19681_ (.A(_03556_),
    .X(_01071_));
 sky130_fd_sc_hd__buf_1 _19682_ (.A(\core.cpuregs[0][17] ),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_1 _19683_ (.A(_03557_),
    .X(_01072_));
 sky130_fd_sc_hd__clkbuf_1 _19684_ (.A(\core.cpuregs[0][18] ),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _19685_ (.A(_03558_),
    .X(_01073_));
 sky130_fd_sc_hd__clkbuf_1 _19686_ (.A(\core.cpuregs[0][19] ),
    .X(_03559_));
 sky130_fd_sc_hd__buf_1 _19687_ (.A(_03559_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_1 _19688_ (.A(\core.cpuregs[0][20] ),
    .X(_03560_));
 sky130_fd_sc_hd__clkbuf_1 _19689_ (.A(_03560_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_1 _19690_ (.A(\core.cpuregs[0][21] ),
    .X(_03561_));
 sky130_fd_sc_hd__buf_1 _19691_ (.A(_03561_),
    .X(_01076_));
 sky130_fd_sc_hd__clkbuf_1 _19692_ (.A(\core.cpuregs[0][22] ),
    .X(_03562_));
 sky130_fd_sc_hd__buf_1 _19693_ (.A(_03562_),
    .X(_01077_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19694_ (.A(\core.cpuregs[0][23] ),
    .X(_03563_));
 sky130_fd_sc_hd__buf_1 _19695_ (.A(_03563_),
    .X(_01078_));
 sky130_fd_sc_hd__clkbuf_1 _19696_ (.A(\core.cpuregs[0][24] ),
    .X(_03564_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19697_ (.A(_03564_),
    .X(_01079_));
 sky130_fd_sc_hd__clkbuf_1 _19698_ (.A(\core.cpuregs[0][25] ),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _19699_ (.A(_03565_),
    .X(_01080_));
 sky130_fd_sc_hd__buf_1 _19700_ (.A(\core.cpuregs[0][26] ),
    .X(_03566_));
 sky130_fd_sc_hd__buf_1 _19701_ (.A(_03566_),
    .X(_01081_));
 sky130_fd_sc_hd__clkbuf_1 _19702_ (.A(\core.cpuregs[0][27] ),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _19703_ (.A(_03567_),
    .X(_01082_));
 sky130_fd_sc_hd__clkbuf_1 _19704_ (.A(\core.cpuregs[0][28] ),
    .X(_03568_));
 sky130_fd_sc_hd__buf_1 _19705_ (.A(_03568_),
    .X(_01083_));
 sky130_fd_sc_hd__clkbuf_1 _19706_ (.A(\core.cpuregs[0][29] ),
    .X(_03569_));
 sky130_fd_sc_hd__buf_1 _19707_ (.A(_03569_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_1 _19708_ (.A(\core.cpuregs[0][30] ),
    .X(_03570_));
 sky130_fd_sc_hd__buf_1 _19709_ (.A(_03570_),
    .X(_01085_));
 sky130_fd_sc_hd__buf_1 _19710_ (.A(\core.cpuregs[0][31] ),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _19711_ (.A(_03571_),
    .X(_01086_));
 sky130_fd_sc_hd__nor2_8 _19712_ (.A(_03396_),
    .B(_09950_),
    .Y(_03572_));
 sky130_fd_sc_hd__clkbuf_2 _19713_ (.A(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_2 _19714_ (.A(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _19715_ (.A0(\core.cpuregs[8][0] ),
    .A1(_03455_),
    .S(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__clkbuf_2 _19716_ (.A(_03575_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_2 _19717_ (.A0(\core.cpuregs[8][1] ),
    .A1(_03459_),
    .S(_03574_),
    .X(_03576_));
 sky130_fd_sc_hd__buf_1 _19718_ (.A(_03576_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_2 _19719_ (.A(_03573_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _19720_ (.A0(\core.cpuregs[8][2] ),
    .A1(_03461_),
    .S(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__buf_1 _19721_ (.A(_03578_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _19722_ (.A0(\core.cpuregs[8][3] ),
    .A1(_03463_),
    .S(_03577_),
    .X(_03579_));
 sky130_fd_sc_hd__buf_1 _19723_ (.A(_03579_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_2 _19724_ (.A0(\core.cpuregs[8][4] ),
    .A1(_03465_),
    .S(_03577_),
    .X(_03580_));
 sky130_fd_sc_hd__buf_1 _19725_ (.A(_03580_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _19726_ (.A0(\core.cpuregs[8][5] ),
    .A1(_03467_),
    .S(_03577_),
    .X(_03581_));
 sky130_fd_sc_hd__clkbuf_1 _19727_ (.A(_03581_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _19728_ (.A0(\core.cpuregs[8][6] ),
    .A1(_03469_),
    .S(_03577_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_1 _19729_ (.A(_03582_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _19730_ (.A0(\core.cpuregs[8][7] ),
    .A1(_03472_),
    .S(_03577_),
    .X(_03583_));
 sky130_fd_sc_hd__buf_1 _19731_ (.A(_03583_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _19732_ (.A0(\core.cpuregs[8][8] ),
    .A1(_03474_),
    .S(_03573_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _19733_ (.A(_03584_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _19734_ (.A0(\core.cpuregs[8][9] ),
    .A1(_03476_),
    .S(_03573_),
    .X(_03585_));
 sky130_fd_sc_hd__buf_1 _19735_ (.A(_03585_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _19736_ (.A0(\core.cpuregs[8][10] ),
    .A1(_03478_),
    .S(_03573_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _19737_ (.A(_03586_),
    .X(_01097_));
 sky130_fd_sc_hd__inv_2 _19738_ (.A(_03572_),
    .Y(_03587_));
 sky130_fd_sc_hd__clkbuf_4 _19739_ (.A(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__mux2_1 _19740_ (.A0(_03480_),
    .A1(\core.cpuregs[8][11] ),
    .S(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__clkbuf_1 _19741_ (.A(_03589_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _19742_ (.A0(\core.cpuregs[8][12] ),
    .A1(_03485_),
    .S(_03573_),
    .X(_03590_));
 sky130_fd_sc_hd__buf_4 _19743_ (.A(_03590_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _19744_ (.A0(_03487_),
    .A1(\core.cpuregs[8][13] ),
    .S(_03588_),
    .X(_03591_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19745_ (.A(_03591_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _19746_ (.A0(_03489_),
    .A1(\core.cpuregs[8][14] ),
    .S(_03587_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _19747_ (.A(_03592_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _19748_ (.A0(_03491_),
    .A1(\core.cpuregs[8][15] ),
    .S(_03587_),
    .X(_03593_));
 sky130_fd_sc_hd__clkbuf_1 _19749_ (.A(_03593_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _19750_ (.A0(_03493_),
    .A1(\core.cpuregs[8][16] ),
    .S(_03587_),
    .X(_03594_));
 sky130_fd_sc_hd__clkbuf_1 _19751_ (.A(_03594_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _19752_ (.A0(_03495_),
    .A1(\core.cpuregs[8][17] ),
    .S(_03587_),
    .X(_03595_));
 sky130_fd_sc_hd__clkbuf_1 _19753_ (.A(_03595_),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_4 _19754_ (.A(_09441_),
    .X(_03596_));
 sky130_fd_sc_hd__and2_1 _19755_ (.A(_03588_),
    .B(\core.cpuregs[8][18] ),
    .X(_03597_));
 sky130_fd_sc_hd__a21o_1 _19756_ (.A1(_03596_),
    .A2(_03574_),
    .B1(_03597_),
    .X(_01105_));
 sky130_fd_sc_hd__clkbuf_4 _19757_ (.A(_03574_),
    .X(_03598_));
 sky130_fd_sc_hd__nand2_1 _19758_ (.A(_03130_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19759_ (.A(_03588_),
    .X(_03600_));
 sky130_fd_sc_hd__nand2_1 _19760_ (.A(_03600_),
    .B(\core.cpuregs[8][19] ),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _19761_ (.A(_03599_),
    .B(_03601_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_1 _19762_ (.A(_03502_),
    .B(_03598_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand2_1 _19763_ (.A(_03600_),
    .B(\core.cpuregs[8][20] ),
    .Y(_03603_));
 sky130_fd_sc_hd__nand2_1 _19764_ (.A(_03602_),
    .B(_03603_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_1 _19765_ (.A(_03508_),
    .B(_03598_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand2_1 _19766_ (.A(_03600_),
    .B(net165),
    .Y(_03605_));
 sky130_fd_sc_hd__nand2_1 _19767_ (.A(_03604_),
    .B(_03605_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand2_1 _19768_ (.A(_03141_),
    .B(_03598_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand2_1 _19769_ (.A(_03600_),
    .B(\core.cpuregs[8][22] ),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_1 _19770_ (.A(_03606_),
    .B(_03607_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _19771_ (.A(_03513_),
    .B(_03598_),
    .Y(_03608_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(_03600_),
    .B(net146),
    .Y(_03609_));
 sky130_fd_sc_hd__nand2_1 _19773_ (.A(_03608_),
    .B(_03609_),
    .Y(_01110_));
 sky130_fd_sc_hd__nand2_2 _19774_ (.A(_03516_),
    .B(_03598_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand2_1 _19775_ (.A(_03600_),
    .B(net149),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _19776_ (.A(_03610_),
    .B(_03611_),
    .Y(_01111_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19777_ (.A(_03574_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _19778_ (.A(_03519_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19779_ (.A(_03588_),
    .X(_03614_));
 sky130_fd_sc_hd__nand2_1 _19780_ (.A(_03614_),
    .B(\core.cpuregs[8][25] ),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_2 _19781_ (.A(_03613_),
    .B(_03615_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _19782_ (.A(_03522_),
    .B(_03612_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_2 _19783_ (.A(_03614_),
    .B(net143),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _19784_ (.A(_03616_),
    .B(_03617_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _19785_ (.A(_03525_),
    .B(_03612_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _19786_ (.A(_03614_),
    .B(\core.cpuregs[8][27] ),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _19787_ (.A(_03618_),
    .B(_03619_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2_2 _19788_ (.A(_03528_),
    .B(_03612_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_1 _19789_ (.A(_03614_),
    .B(\core.cpuregs[8][28] ),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_1 _19790_ (.A(_03620_),
    .B(_03621_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _19791_ (.A(_03531_),
    .B(_03612_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2_1 _19792_ (.A(_03614_),
    .B(\core.cpuregs[8][29] ),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _19793_ (.A(_03622_),
    .B(_03623_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _19794_ (.A(_03534_),
    .B(_03612_),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _19795_ (.A(_03614_),
    .B(net155),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _19796_ (.A(_03624_),
    .B(_03625_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _19797_ (.A(_03537_),
    .B(_03574_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _19798_ (.A(_03588_),
    .B(\core.cpuregs[8][31] ),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _19799_ (.A(_03626_),
    .B(_03627_),
    .Y(_01118_));
 sky130_fd_sc_hd__and3_1 _19800_ (.A(_09317_),
    .B(_09318_),
    .C(\core.latched_rd[2] ),
    .X(_03628_));
 sky130_fd_sc_hd__inv_2 _19801_ (.A(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_1 _19802_ (.A(_03629_),
    .B(_09812_),
    .Y(_03630_));
 sky130_fd_sc_hd__clkbuf_2 _19803_ (.A(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _19804_ (.A0(\core.cpuregs[7][0] ),
    .A1(_03455_),
    .S(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _19805_ (.A(_03632_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _19806_ (.A0(\core.cpuregs[7][1] ),
    .A1(_03459_),
    .S(_03631_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_1 _19807_ (.A(_03633_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _19808_ (.A0(\core.cpuregs[7][2] ),
    .A1(_03461_),
    .S(_03631_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _19809_ (.A(_03634_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _19810_ (.A0(\core.cpuregs[7][3] ),
    .A1(_03463_),
    .S(_03631_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _19811_ (.A(_03635_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _19812_ (.A0(\core.cpuregs[7][4] ),
    .A1(_03465_),
    .S(_03631_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _19813_ (.A(_03636_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _19814_ (.A0(\core.cpuregs[7][5] ),
    .A1(_03467_),
    .S(_03631_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _19815_ (.A(_03637_),
    .X(_01124_));
 sky130_fd_sc_hd__clkbuf_4 _19816_ (.A(_03630_),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _19817_ (.A0(\core.cpuregs[7][6] ),
    .A1(_03469_),
    .S(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_1 _19818_ (.A(_03639_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_2 _19819_ (.A0(\core.cpuregs[7][7] ),
    .A1(_03472_),
    .S(_03638_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_1 _19820_ (.A(_03640_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _19821_ (.A0(\core.cpuregs[7][8] ),
    .A1(_03474_),
    .S(_03638_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _19822_ (.A(_03641_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _19823_ (.A0(\core.cpuregs[7][9] ),
    .A1(_03476_),
    .S(_03638_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_1 _19824_ (.A(_03642_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _19825_ (.A0(\core.cpuregs[7][10] ),
    .A1(_03478_),
    .S(_03638_),
    .X(_03643_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19826_ (.A(_03643_),
    .X(_01129_));
 sky130_fd_sc_hd__and3_1 _19827_ (.A(_09324_),
    .B(_09326_),
    .C(_03628_),
    .X(_03644_));
 sky130_fd_sc_hd__inv_2 _19828_ (.A(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__clkbuf_4 _19829_ (.A(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _19830_ (.A0(_03480_),
    .A1(\core.cpuregs[7][11] ),
    .S(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _19831_ (.A(_03647_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _19832_ (.A0(\core.cpuregs[7][12] ),
    .A1(_03485_),
    .S(_03638_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_4 _19833_ (.A(_03648_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _19834_ (.A0(_03487_),
    .A1(\core.cpuregs[7][13] ),
    .S(_03646_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _19835_ (.A(_03649_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _19836_ (.A0(_03489_),
    .A1(\core.cpuregs[7][14] ),
    .S(_03646_),
    .X(_03650_));
 sky130_fd_sc_hd__clkbuf_1 _19837_ (.A(_03650_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _19838_ (.A0(_03491_),
    .A1(\core.cpuregs[7][15] ),
    .S(_03646_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _19839_ (.A(_03651_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _19840_ (.A0(_03493_),
    .A1(\core.cpuregs[7][16] ),
    .S(_03646_),
    .X(_03652_));
 sky130_fd_sc_hd__clkbuf_1 _19841_ (.A(_03652_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _19842_ (.A0(_03495_),
    .A1(\core.cpuregs[7][17] ),
    .S(_03645_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_1 _19843_ (.A(_03653_),
    .X(_01136_));
 sky130_fd_sc_hd__buf_4 _19844_ (.A(_03630_),
    .X(_03654_));
 sky130_fd_sc_hd__and2_1 _19845_ (.A(_03646_),
    .B(\core.cpuregs[7][18] ),
    .X(_03655_));
 sky130_fd_sc_hd__a21o_1 _19846_ (.A1(_03596_),
    .A2(_03654_),
    .B1(_03655_),
    .X(_01137_));
 sky130_fd_sc_hd__inv_2 _19847_ (.A(\core.cpuregs[7][19] ),
    .Y(_03656_));
 sky130_fd_sc_hd__clkbuf_4 _19848_ (.A(_03654_),
    .X(_03657_));
 sky130_fd_sc_hd__nand2_1 _19849_ (.A(_09447_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_2 _19850_ (.A1(_03656_),
    .A2(_03654_),
    .B1(_03658_),
    .Y(_01138_));
 sky130_fd_sc_hd__buf_4 _19851_ (.A(_03654_),
    .X(_03659_));
 sky130_fd_sc_hd__nand2_4 _19852_ (.A(_03502_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19853_ (.A(_03645_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_4 _19854_ (.A(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__nand2_1 _19855_ (.A(_03662_),
    .B(\core.cpuregs[7][20] ),
    .Y(_03663_));
 sky130_fd_sc_hd__nand2_2 _19856_ (.A(_03660_),
    .B(_03663_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _19857_ (.A(_03508_),
    .B(_03659_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_2 _19858_ (.A(_03662_),
    .B(\core.cpuregs[7][21] ),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _19859_ (.A(_03664_),
    .B(_03665_),
    .Y(_01140_));
 sky130_fd_sc_hd__inv_2 _19860_ (.A(\core.cpuregs[7][22] ),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _19861_ (.A(_09473_),
    .B(_03654_),
    .Y(_03667_));
 sky130_fd_sc_hd__o21ai_2 _19862_ (.A1(_03666_),
    .A2(_03654_),
    .B1(_03667_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand2_1 _19863_ (.A(_03513_),
    .B(_03659_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand2_1 _19864_ (.A(_03662_),
    .B(net126),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _19865_ (.A(_03668_),
    .B(_03669_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_1 _19866_ (.A(_03516_),
    .B(_03659_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _19867_ (.A(_03662_),
    .B(\core.cpuregs[7][24] ),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _19868_ (.A(_03670_),
    .B(_03671_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand2_1 _19869_ (.A(_03519_),
    .B(_03659_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _19870_ (.A(_03662_),
    .B(\core.cpuregs[7][25] ),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _19871_ (.A(_03672_),
    .B(_03673_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_1 _19872_ (.A(_03522_),
    .B(_03659_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _19873_ (.A(_03662_),
    .B(net187),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _19874_ (.A(_03674_),
    .B(_03675_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _19875_ (.A(_03525_),
    .B(_03657_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand2_1 _19876_ (.A(_03661_),
    .B(\core.cpuregs[7][27] ),
    .Y(_03677_));
 sky130_fd_sc_hd__nand2_2 _19877_ (.A(_03676_),
    .B(_03677_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand2_2 _19878_ (.A(_03528_),
    .B(_03657_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand2_1 _19879_ (.A(_03661_),
    .B(\core.cpuregs[7][28] ),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_1 _19880_ (.A(_03678_),
    .B(_03679_),
    .Y(_01147_));
 sky130_fd_sc_hd__nand2_1 _19881_ (.A(_03531_),
    .B(_03657_),
    .Y(_03680_));
 sky130_fd_sc_hd__nand2_1 _19882_ (.A(_03661_),
    .B(\core.cpuregs[7][29] ),
    .Y(_03681_));
 sky130_fd_sc_hd__nand2_1 _19883_ (.A(_03680_),
    .B(_03681_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2_1 _19884_ (.A(_03534_),
    .B(_03657_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _19885_ (.A(_03661_),
    .B(\core.cpuregs[7][30] ),
    .Y(_03683_));
 sky130_fd_sc_hd__nand2_1 _19886_ (.A(_03682_),
    .B(_03683_),
    .Y(_01149_));
 sky130_fd_sc_hd__nand2_1 _19887_ (.A(_03537_),
    .B(_03657_),
    .Y(_03684_));
 sky130_fd_sc_hd__nand2_1 _19888_ (.A(_03661_),
    .B(\core.cpuregs[7][31] ),
    .Y(_03685_));
 sky130_fd_sc_hd__nand2_1 _19889_ (.A(_03684_),
    .B(_03685_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _19890_ (.A(_03629_),
    .B(_10158_),
    .Y(_03686_));
 sky130_fd_sc_hd__clkbuf_4 _19891_ (.A(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_2 _19892_ (.A(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_2 _19893_ (.A0(\core.cpuregs[6][0] ),
    .A1(_03455_),
    .S(_03688_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _19894_ (.A(_03689_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _19895_ (.A0(\core.cpuregs[6][1] ),
    .A1(_03459_),
    .S(_03688_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _19896_ (.A(_03690_),
    .X(_01152_));
 sky130_fd_sc_hd__clkbuf_4 _19897_ (.A(_03687_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _19898_ (.A0(\core.cpuregs[6][2] ),
    .A1(_03461_),
    .S(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__buf_1 _19899_ (.A(_03692_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(\core.cpuregs[6][3] ),
    .A1(_03463_),
    .S(_03691_),
    .X(_03693_));
 sky130_fd_sc_hd__buf_1 _19901_ (.A(_03693_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _19902_ (.A0(\core.cpuregs[6][4] ),
    .A1(_03465_),
    .S(_03691_),
    .X(_03694_));
 sky130_fd_sc_hd__clkbuf_1 _19903_ (.A(_03694_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _19904_ (.A0(\core.cpuregs[6][5] ),
    .A1(_03467_),
    .S(_03691_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_1 _19905_ (.A(_03695_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _19906_ (.A0(\core.cpuregs[6][6] ),
    .A1(_03469_),
    .S(_03691_),
    .X(_03696_));
 sky130_fd_sc_hd__buf_4 _19907_ (.A(_03696_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _19908_ (.A0(\core.cpuregs[6][7] ),
    .A1(_03472_),
    .S(_03691_),
    .X(_03697_));
 sky130_fd_sc_hd__buf_4 _19909_ (.A(_03697_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _19910_ (.A0(\core.cpuregs[6][8] ),
    .A1(_03474_),
    .S(_03687_),
    .X(_03698_));
 sky130_fd_sc_hd__buf_1 _19911_ (.A(_03698_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _19912_ (.A0(\core.cpuregs[6][9] ),
    .A1(_03476_),
    .S(_03687_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_1 _19913_ (.A(_03699_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _19914_ (.A0(\core.cpuregs[6][10] ),
    .A1(_03478_),
    .S(_03687_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_1 _19915_ (.A(_03700_),
    .X(_01161_));
 sky130_fd_sc_hd__inv_2 _19916_ (.A(_03686_),
    .Y(_03701_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19917_ (.A(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _19918_ (.A0(_03480_),
    .A1(\core.cpuregs[6][11] ),
    .S(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_1 _19919_ (.A(_03703_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _19920_ (.A0(\core.cpuregs[6][12] ),
    .A1(_03485_),
    .S(_03687_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_1 _19921_ (.A(_03704_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _19922_ (.A0(_03487_),
    .A1(\core.cpuregs[6][13] ),
    .S(_03702_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_1 _19923_ (.A(_03705_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_2 _19924_ (.A0(_03489_),
    .A1(\core.cpuregs[6][14] ),
    .S(_03701_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_2 _19925_ (.A(_03706_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _19926_ (.A0(_03491_),
    .A1(\core.cpuregs[6][15] ),
    .S(_03701_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_1 _19927_ (.A(_03707_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _19928_ (.A0(_03493_),
    .A1(\core.cpuregs[6][16] ),
    .S(_03701_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _19929_ (.A(_03708_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _19930_ (.A0(_03495_),
    .A1(\core.cpuregs[6][17] ),
    .S(_03701_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_1 _19931_ (.A(_03709_),
    .X(_01168_));
 sky130_fd_sc_hd__and2_1 _19932_ (.A(_03702_),
    .B(\core.cpuregs[6][18] ),
    .X(_03710_));
 sky130_fd_sc_hd__a21o_1 _19933_ (.A1(_03596_),
    .A2(_03688_),
    .B1(_03710_),
    .X(_01169_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19934_ (.A(_09447_),
    .X(_03711_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19935_ (.A(_03688_),
    .X(_03712_));
 sky130_fd_sc_hd__nand2_1 _19936_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__clkbuf_2 _19937_ (.A(_03702_),
    .X(_03714_));
 sky130_fd_sc_hd__nand2_1 _19938_ (.A(_03714_),
    .B(\core.cpuregs[6][19] ),
    .Y(_03715_));
 sky130_fd_sc_hd__nand2_1 _19939_ (.A(_03713_),
    .B(_03715_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_2 _19940_ (.A(_03502_),
    .B(_03712_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _19941_ (.A(_03714_),
    .B(\core.cpuregs[6][20] ),
    .Y(_03717_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(_03716_),
    .B(_03717_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _19943_ (.A(_03508_),
    .B(_03712_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_2 _19944_ (.A(_03714_),
    .B(\core.cpuregs[6][21] ),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _19945_ (.A(_03718_),
    .B(_03719_),
    .Y(_01172_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19946_ (.A(_09473_),
    .X(_03720_));
 sky130_fd_sc_hd__nand2_1 _19947_ (.A(_03720_),
    .B(_03712_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _19948_ (.A(_03714_),
    .B(\core.cpuregs[6][22] ),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _19949_ (.A(_03721_),
    .B(_03722_),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _19950_ (.A(_03513_),
    .B(_03712_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand2_1 _19951_ (.A(_03714_),
    .B(\core.cpuregs[6][23] ),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_1 _19952_ (.A(_03723_),
    .B(_03724_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(_03516_),
    .B(_03712_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_2 _19954_ (.A(_03714_),
    .B(\core.cpuregs[6][24] ),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2_1 _19955_ (.A(_03725_),
    .B(_03726_),
    .Y(_01175_));
 sky130_fd_sc_hd__clkbuf_2 _19956_ (.A(_03688_),
    .X(_03727_));
 sky130_fd_sc_hd__nand2_1 _19957_ (.A(_03519_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__buf_4 _19958_ (.A(_03702_),
    .X(_03729_));
 sky130_fd_sc_hd__nand2_1 _19959_ (.A(_03729_),
    .B(net197),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _19960_ (.A(_03728_),
    .B(_03730_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_2 _19961_ (.A(_03522_),
    .B(_03727_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _19962_ (.A(_03729_),
    .B(\core.cpuregs[6][26] ),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_2 _19963_ (.A(_03731_),
    .B(_03732_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_1 _19964_ (.A(_03525_),
    .B(_03727_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2_1 _19965_ (.A(_03729_),
    .B(\core.cpuregs[6][27] ),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _19966_ (.A(_03733_),
    .B(_03734_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_2 _19967_ (.A(_03528_),
    .B(_03727_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_1 _19968_ (.A(_03729_),
    .B(\core.cpuregs[6][28] ),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _19969_ (.A(_03735_),
    .B(_03736_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _19970_ (.A(_03531_),
    .B(_03727_),
    .Y(_03737_));
 sky130_fd_sc_hd__nand2_2 _19971_ (.A(_03729_),
    .B(\core.cpuregs[6][29] ),
    .Y(_03738_));
 sky130_fd_sc_hd__nand2_1 _19972_ (.A(_03737_),
    .B(_03738_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _19973_ (.A(_03534_),
    .B(_03727_),
    .Y(_03739_));
 sky130_fd_sc_hd__nand2_1 _19974_ (.A(_03729_),
    .B(net151),
    .Y(_03740_));
 sky130_fd_sc_hd__nand2_1 _19975_ (.A(_03739_),
    .B(_03740_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _19976_ (.A(_03537_),
    .B(_03688_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _19977_ (.A(_03702_),
    .B(net134),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _19978_ (.A(_03741_),
    .B(_03742_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _19979_ (.A(_03629_),
    .B(_02778_),
    .Y(_03743_));
 sky130_fd_sc_hd__clkbuf_2 _19980_ (.A(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_2 _19981_ (.A(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _19982_ (.A0(\core.cpuregs[5][0] ),
    .A1(_03455_),
    .S(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _19983_ (.A(_03746_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _19984_ (.A0(\core.cpuregs[5][1] ),
    .A1(_03459_),
    .S(_03745_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _19985_ (.A(_03747_),
    .X(_01184_));
 sky130_fd_sc_hd__buf_2 _19986_ (.A(_03744_),
    .X(_03748_));
 sky130_fd_sc_hd__mux2_1 _19987_ (.A0(\core.cpuregs[5][2] ),
    .A1(_03461_),
    .S(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _19988_ (.A(_03749_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _19989_ (.A0(\core.cpuregs[5][3] ),
    .A1(_03463_),
    .S(_03748_),
    .X(_03750_));
 sky130_fd_sc_hd__buf_1 _19990_ (.A(_03750_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _19991_ (.A0(\core.cpuregs[5][4] ),
    .A1(_03465_),
    .S(_03748_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _19992_ (.A(_03751_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _19993_ (.A0(\core.cpuregs[5][5] ),
    .A1(_03467_),
    .S(_03748_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _19994_ (.A(_03752_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _19995_ (.A0(\core.cpuregs[5][6] ),
    .A1(_03469_),
    .S(_03748_),
    .X(_03753_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19996_ (.A(_03753_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _19997_ (.A0(\core.cpuregs[5][7] ),
    .A1(_03472_),
    .S(_03748_),
    .X(_03754_));
 sky130_fd_sc_hd__buf_1 _19998_ (.A(_03754_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _19999_ (.A0(\core.cpuregs[5][8] ),
    .A1(_03474_),
    .S(_03744_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _20000_ (.A(_03755_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _20001_ (.A0(\core.cpuregs[5][9] ),
    .A1(_03476_),
    .S(_03744_),
    .X(_03756_));
 sky130_fd_sc_hd__buf_4 _20002_ (.A(_03756_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _20003_ (.A0(\core.cpuregs[5][10] ),
    .A1(_03478_),
    .S(_03744_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _20004_ (.A(_03757_),
    .X(_01193_));
 sky130_fd_sc_hd__inv_2 _20005_ (.A(_03743_),
    .Y(_03758_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20006_ (.A(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__mux2_1 _20007_ (.A0(_03480_),
    .A1(\core.cpuregs[5][11] ),
    .S(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_4 _20008_ (.A(_03760_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_4 _20009_ (.A0(\core.cpuregs[5][12] ),
    .A1(_03485_),
    .S(_03744_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _20010_ (.A(_03761_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _20011_ (.A0(_03487_),
    .A1(\core.cpuregs[5][13] ),
    .S(_03759_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _20012_ (.A(_03762_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _20013_ (.A0(_03489_),
    .A1(\core.cpuregs[5][14] ),
    .S(_03758_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _20014_ (.A(_03763_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _20015_ (.A0(_03491_),
    .A1(\core.cpuregs[5][15] ),
    .S(_03758_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _20016_ (.A(_03764_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_4 _20017_ (.A0(_03493_),
    .A1(\core.cpuregs[5][16] ),
    .S(_03758_),
    .X(_03765_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20018_ (.A(_03765_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _20019_ (.A0(_03495_),
    .A1(\core.cpuregs[5][17] ),
    .S(_03758_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _20020_ (.A(_03766_),
    .X(_01200_));
 sky130_fd_sc_hd__and2_1 _20021_ (.A(_03759_),
    .B(\core.cpuregs[5][18] ),
    .X(_03767_));
 sky130_fd_sc_hd__a21o_1 _20022_ (.A1(_03596_),
    .A2(_03745_),
    .B1(_03767_),
    .X(_01201_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20023_ (.A(_03745_),
    .X(_03768_));
 sky130_fd_sc_hd__nand2_1 _20024_ (.A(_03711_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__clkbuf_4 _20025_ (.A(_03759_),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_1 _20026_ (.A(_03770_),
    .B(\core.cpuregs[5][19] ),
    .Y(_03771_));
 sky130_fd_sc_hd__nand2_1 _20027_ (.A(_03769_),
    .B(_03771_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _20028_ (.A(_03502_),
    .B(_03768_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _20029_ (.A(_03770_),
    .B(\core.cpuregs[5][20] ),
    .Y(_03773_));
 sky130_fd_sc_hd__nand2_1 _20030_ (.A(_03772_),
    .B(_03773_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _20031_ (.A(_03508_),
    .B(_03768_),
    .Y(_03774_));
 sky130_fd_sc_hd__nand2_1 _20032_ (.A(_03770_),
    .B(\core.cpuregs[5][21] ),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _20033_ (.A(_03774_),
    .B(_03775_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _20034_ (.A(_03720_),
    .B(_03768_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand2_2 _20035_ (.A(_03770_),
    .B(\core.cpuregs[5][22] ),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _20036_ (.A(_03776_),
    .B(_03777_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _20037_ (.A(_03513_),
    .B(_03768_),
    .Y(_03778_));
 sky130_fd_sc_hd__nand2_1 _20038_ (.A(_03770_),
    .B(net163),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2_1 _20039_ (.A(_03778_),
    .B(_03779_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _20040_ (.A(_03516_),
    .B(_03768_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _20041_ (.A(_03770_),
    .B(\core.cpuregs[5][24] ),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_1 _20042_ (.A(_03780_),
    .B(_03781_),
    .Y(_01207_));
 sky130_fd_sc_hd__buf_2 _20043_ (.A(_03745_),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _20044_ (.A(_03519_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20045_ (.A(_03759_),
    .X(_03784_));
 sky130_fd_sc_hd__nand2_1 _20046_ (.A(_03784_),
    .B(\core.cpuregs[5][25] ),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2_1 _20047_ (.A(_03783_),
    .B(_03785_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_1 _20048_ (.A(_03522_),
    .B(_03782_),
    .Y(_03786_));
 sky130_fd_sc_hd__nand2_1 _20049_ (.A(_03784_),
    .B(\core.cpuregs[5][26] ),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _20050_ (.A(_03786_),
    .B(_03787_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_2 _20051_ (.A(_03525_),
    .B(_03782_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _20052_ (.A(_03784_),
    .B(\core.cpuregs[5][27] ),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _20053_ (.A(_03788_),
    .B(_03789_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_2 _20054_ (.A(_03528_),
    .B(_03782_),
    .Y(_03790_));
 sky130_fd_sc_hd__nand2_1 _20055_ (.A(_03784_),
    .B(\core.cpuregs[5][28] ),
    .Y(_03791_));
 sky130_fd_sc_hd__nand2_1 _20056_ (.A(_03790_),
    .B(_03791_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _20057_ (.A(_03531_),
    .B(_03782_),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2_1 _20058_ (.A(_03784_),
    .B(\core.cpuregs[5][29] ),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _20059_ (.A(_03792_),
    .B(_03793_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_1 _20060_ (.A(_03534_),
    .B(_03782_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_1 _20061_ (.A(_03784_),
    .B(\core.cpuregs[5][30] ),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _20062_ (.A(_03794_),
    .B(_03795_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand2_1 _20063_ (.A(_03537_),
    .B(_03745_),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _20064_ (.A(_03759_),
    .B(net178),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _20065_ (.A(_03796_),
    .B(_03797_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _20066_ (.A(_03629_),
    .B(_09950_),
    .Y(_03798_));
 sky130_fd_sc_hd__buf_4 _20067_ (.A(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__clkbuf_2 _20068_ (.A(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_1 _20069_ (.A0(\core.cpuregs[4][0] ),
    .A1(_03455_),
    .S(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__clkbuf_1 _20070_ (.A(_03801_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _20071_ (.A0(\core.cpuregs[4][1] ),
    .A1(_03459_),
    .S(_03800_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _20072_ (.A(_03802_),
    .X(_01216_));
 sky130_fd_sc_hd__clkbuf_2 _20073_ (.A(_03799_),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_1 _20074_ (.A0(\core.cpuregs[4][2] ),
    .A1(_03461_),
    .S(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _20075_ (.A(_03804_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _20076_ (.A0(\core.cpuregs[4][3] ),
    .A1(_03463_),
    .S(_03803_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _20077_ (.A(_03805_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _20078_ (.A0(\core.cpuregs[4][4] ),
    .A1(_03465_),
    .S(_03803_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _20079_ (.A(_03806_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _20080_ (.A0(\core.cpuregs[4][5] ),
    .A1(_03467_),
    .S(_03803_),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_1 _20081_ (.A(_03807_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _20082_ (.A0(\core.cpuregs[4][6] ),
    .A1(_03469_),
    .S(_03803_),
    .X(_03808_));
 sky130_fd_sc_hd__buf_1 _20083_ (.A(_03808_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_4 _20084_ (.A0(\core.cpuregs[4][7] ),
    .A1(_03472_),
    .S(_03803_),
    .X(_03809_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20085_ (.A(_03809_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _20086_ (.A0(\core.cpuregs[4][8] ),
    .A1(_03474_),
    .S(_03799_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _20087_ (.A(_03810_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _20088_ (.A0(\core.cpuregs[4][9] ),
    .A1(_03476_),
    .S(_03799_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _20089_ (.A(_03811_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _20090_ (.A0(\core.cpuregs[4][10] ),
    .A1(_03478_),
    .S(_03799_),
    .X(_03812_));
 sky130_fd_sc_hd__buf_1 _20091_ (.A(_03812_),
    .X(_01225_));
 sky130_fd_sc_hd__inv_2 _20092_ (.A(_03798_),
    .Y(_03813_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20093_ (.A(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__mux2_1 _20094_ (.A0(_03480_),
    .A1(\core.cpuregs[4][11] ),
    .S(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _20095_ (.A(_03815_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _20096_ (.A0(\core.cpuregs[4][12] ),
    .A1(_03485_),
    .S(_03799_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _20097_ (.A(_03816_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _20098_ (.A0(_03487_),
    .A1(\core.cpuregs[4][13] ),
    .S(_03814_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _20099_ (.A(_03817_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _20100_ (.A0(_03489_),
    .A1(\core.cpuregs[4][14] ),
    .S(_03813_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _20101_ (.A(_03818_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _20102_ (.A0(_03491_),
    .A1(\core.cpuregs[4][15] ),
    .S(_03813_),
    .X(_03819_));
 sky130_fd_sc_hd__clkbuf_1 _20103_ (.A(_03819_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_2 _20104_ (.A0(_03493_),
    .A1(\core.cpuregs[4][16] ),
    .S(_03813_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_8 _20105_ (.A(_03820_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _20106_ (.A0(_03495_),
    .A1(\core.cpuregs[4][17] ),
    .S(_03813_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _20107_ (.A(_03821_),
    .X(_01232_));
 sky130_fd_sc_hd__and2_1 _20108_ (.A(_03814_),
    .B(\core.cpuregs[4][18] ),
    .X(_03822_));
 sky130_fd_sc_hd__a21o_1 _20109_ (.A1(_03596_),
    .A2(_03800_),
    .B1(_03822_),
    .X(_01233_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20110_ (.A(_03800_),
    .X(_03823_));
 sky130_fd_sc_hd__nand2_1 _20111_ (.A(_03711_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20112_ (.A(_03814_),
    .X(_03825_));
 sky130_fd_sc_hd__nand2_1 _20113_ (.A(_03825_),
    .B(\core.cpuregs[4][19] ),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_03824_),
    .B(_03826_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand2_1 _20115_ (.A(_03502_),
    .B(_03823_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _20116_ (.A(_03825_),
    .B(\core.cpuregs[4][20] ),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _20117_ (.A(_03827_),
    .B(_03828_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_1 _20118_ (.A(_03508_),
    .B(_03823_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_1 _20119_ (.A(_03825_),
    .B(\core.cpuregs[4][21] ),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _20120_ (.A(_03829_),
    .B(_03830_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(_03720_),
    .B(_03823_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _20122_ (.A(_03825_),
    .B(net186),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _20123_ (.A(_03831_),
    .B(_03832_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _20124_ (.A(_03513_),
    .B(_03823_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _20125_ (.A(_03825_),
    .B(net172),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_2 _20126_ (.A(_03833_),
    .B(_03834_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _20127_ (.A(_03516_),
    .B(_03823_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_1 _20128_ (.A(_03825_),
    .B(net166),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _20129_ (.A(_03835_),
    .B(_03836_),
    .Y(_01239_));
 sky130_fd_sc_hd__clkbuf_4 _20130_ (.A(_03800_),
    .X(_03837_));
 sky130_fd_sc_hd__nand2_1 _20131_ (.A(_03519_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20132_ (.A(_03814_),
    .X(_03839_));
 sky130_fd_sc_hd__nand2_1 _20133_ (.A(_03839_),
    .B(\core.cpuregs[4][25] ),
    .Y(_03840_));
 sky130_fd_sc_hd__nand2_1 _20134_ (.A(_03838_),
    .B(_03840_),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _20135_ (.A(_03522_),
    .B(_03837_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _20136_ (.A(_03839_),
    .B(\core.cpuregs[4][26] ),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _20137_ (.A(_03841_),
    .B(_03842_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _20138_ (.A(_03525_),
    .B(_03837_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _20139_ (.A(_03839_),
    .B(\core.cpuregs[4][27] ),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _20140_ (.A(_03843_),
    .B(_03844_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_2 _20141_ (.A(_03528_),
    .B(_03837_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _20142_ (.A(_03839_),
    .B(\core.cpuregs[4][28] ),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_2 _20143_ (.A(_03845_),
    .B(_03846_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_2 _20144_ (.A(_03531_),
    .B(_03837_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand2_1 _20145_ (.A(_03839_),
    .B(\core.cpuregs[4][29] ),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2_1 _20146_ (.A(_03847_),
    .B(_03848_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2_1 _20147_ (.A(_03534_),
    .B(_03837_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2_1 _20148_ (.A(_03839_),
    .B(\core.cpuregs[4][30] ),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _20149_ (.A(_03849_),
    .B(_03850_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _20150_ (.A(_03537_),
    .B(_03800_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _20151_ (.A(_03814_),
    .B(net157),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _20152_ (.A(_03851_),
    .B(_03852_),
    .Y(_01246_));
 sky130_fd_sc_hd__buf_1 _20153_ (.A(_09314_),
    .X(_03853_));
 sky130_fd_sc_hd__and3_1 _20154_ (.A(_09554_),
    .B(_09326_),
    .C(_09320_),
    .X(_03854_));
 sky130_fd_sc_hd__clkbuf_2 _20155_ (.A(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_2 _20156_ (.A(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _20157_ (.A0(\core.cpuregs[3][0] ),
    .A1(_03853_),
    .S(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__buf_1 _20158_ (.A(_03857_),
    .X(_01247_));
 sky130_fd_sc_hd__buf_1 _20159_ (.A(_09336_),
    .X(_03858_));
 sky130_fd_sc_hd__mux2_1 _20160_ (.A0(\core.cpuregs[3][1] ),
    .A1(_03858_),
    .S(_03856_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_1 _20161_ (.A(_03859_),
    .X(_01248_));
 sky130_fd_sc_hd__buf_2 _20162_ (.A(_09339_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_2 _20163_ (.A(_03855_),
    .X(_03861_));
 sky130_fd_sc_hd__mux2_1 _20164_ (.A0(\core.cpuregs[3][2] ),
    .A1(_03860_),
    .S(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__buf_2 _20165_ (.A(_03862_),
    .X(_01249_));
 sky130_fd_sc_hd__clkbuf_2 _20166_ (.A(_09348_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _20167_ (.A0(\core.cpuregs[3][3] ),
    .A1(_03863_),
    .S(_03861_),
    .X(_03864_));
 sky130_fd_sc_hd__buf_1 _20168_ (.A(_03864_),
    .X(_01250_));
 sky130_fd_sc_hd__buf_2 _20169_ (.A(_09356_),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _20170_ (.A0(\core.cpuregs[3][4] ),
    .A1(_03865_),
    .S(_03861_),
    .X(_03866_));
 sky130_fd_sc_hd__buf_1 _20171_ (.A(_03866_),
    .X(_01251_));
 sky130_fd_sc_hd__buf_2 _20172_ (.A(_09362_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _20173_ (.A0(\core.cpuregs[3][5] ),
    .A1(_03867_),
    .S(_03861_),
    .X(_03868_));
 sky130_fd_sc_hd__buf_1 _20174_ (.A(_03868_),
    .X(_01252_));
 sky130_fd_sc_hd__buf_2 _20175_ (.A(_09368_),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_1 _20176_ (.A0(\core.cpuregs[3][6] ),
    .A1(_03869_),
    .S(_03861_),
    .X(_03870_));
 sky130_fd_sc_hd__buf_1 _20177_ (.A(_03870_),
    .X(_01253_));
 sky130_fd_sc_hd__buf_1 _20178_ (.A(_09374_),
    .X(_03871_));
 sky130_fd_sc_hd__mux2_2 _20179_ (.A0(\core.cpuregs[3][7] ),
    .A1(_03871_),
    .S(_03861_),
    .X(_03872_));
 sky130_fd_sc_hd__buf_1 _20180_ (.A(_03872_),
    .X(_01254_));
 sky130_fd_sc_hd__buf_1 _20181_ (.A(_09380_),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _20182_ (.A0(\core.cpuregs[3][8] ),
    .A1(_03873_),
    .S(_03855_),
    .X(_03874_));
 sky130_fd_sc_hd__buf_1 _20183_ (.A(_03874_),
    .X(_01255_));
 sky130_fd_sc_hd__buf_1 _20184_ (.A(_09387_),
    .X(_03875_));
 sky130_fd_sc_hd__mux2_2 _20185_ (.A0(\core.cpuregs[3][9] ),
    .A1(_03875_),
    .S(_03855_),
    .X(_03876_));
 sky130_fd_sc_hd__clkbuf_1 _20186_ (.A(_03876_),
    .X(_01256_));
 sky130_fd_sc_hd__buf_1 _20187_ (.A(_09394_),
    .X(_03877_));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(\core.cpuregs[3][10] ),
    .A1(_03877_),
    .S(_03855_),
    .X(_03878_));
 sky130_fd_sc_hd__clkbuf_1 _20189_ (.A(_03878_),
    .X(_01257_));
 sky130_fd_sc_hd__buf_1 _20190_ (.A(_09400_),
    .X(_03879_));
 sky130_fd_sc_hd__inv_2 _20191_ (.A(_03854_),
    .Y(_03880_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20192_ (.A(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_1 _20193_ (.A0(_03879_),
    .A1(\core.cpuregs[3][11] ),
    .S(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__buf_1 _20194_ (.A(_03882_),
    .X(_01258_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20195_ (.A(_09407_),
    .X(_03883_));
 sky130_fd_sc_hd__mux2_1 _20196_ (.A0(\core.cpuregs[3][12] ),
    .A1(_03883_),
    .S(_03855_),
    .X(_03884_));
 sky130_fd_sc_hd__buf_1 _20197_ (.A(_03884_),
    .X(_01259_));
 sky130_fd_sc_hd__buf_4 _20198_ (.A(_09413_),
    .X(_03885_));
 sky130_fd_sc_hd__mux2_1 _20199_ (.A0(_03885_),
    .A1(\core.cpuregs[3][13] ),
    .S(_03881_),
    .X(_03886_));
 sky130_fd_sc_hd__clkbuf_1 _20200_ (.A(_03886_),
    .X(_01260_));
 sky130_fd_sc_hd__buf_1 _20201_ (.A(_09418_),
    .X(_03887_));
 sky130_fd_sc_hd__mux2_1 _20202_ (.A0(_03887_),
    .A1(\core.cpuregs[3][14] ),
    .S(_03880_),
    .X(_03888_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20203_ (.A(_03888_),
    .X(_01261_));
 sky130_fd_sc_hd__buf_1 _20204_ (.A(_09423_),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_2 _20205_ (.A0(_03889_),
    .A1(\core.cpuregs[3][15] ),
    .S(_03880_),
    .X(_03890_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20206_ (.A(_03890_),
    .X(_01262_));
 sky130_fd_sc_hd__clkbuf_8 _20207_ (.A(_09430_),
    .X(_03891_));
 sky130_fd_sc_hd__mux2_1 _20208_ (.A0(_03891_),
    .A1(\core.cpuregs[3][16] ),
    .S(_03880_),
    .X(_03892_));
 sky130_fd_sc_hd__clkbuf_1 _20209_ (.A(_03892_),
    .X(_01263_));
 sky130_fd_sc_hd__buf_1 _20210_ (.A(_09435_),
    .X(_03893_));
 sky130_fd_sc_hd__mux2_1 _20211_ (.A0(_03893_),
    .A1(\core.cpuregs[3][17] ),
    .S(_03880_),
    .X(_03894_));
 sky130_fd_sc_hd__clkbuf_2 _20212_ (.A(_03894_),
    .X(_01264_));
 sky130_fd_sc_hd__and2_1 _20213_ (.A(_03881_),
    .B(\core.cpuregs[3][18] ),
    .X(_03895_));
 sky130_fd_sc_hd__a21o_1 _20214_ (.A1(_03596_),
    .A2(_03856_),
    .B1(_03895_),
    .X(_01265_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20215_ (.A(_03856_),
    .X(_03896_));
 sky130_fd_sc_hd__nand2_1 _20216_ (.A(_03711_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__clkbuf_2 _20217_ (.A(_03881_),
    .X(_03898_));
 sky130_fd_sc_hd__nand2_1 _20218_ (.A(_03898_),
    .B(\core.cpuregs[3][19] ),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _20219_ (.A(_03897_),
    .B(_03899_),
    .Y(_01266_));
 sky130_fd_sc_hd__clkbuf_2 _20220_ (.A(_09457_),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_2 _20221_ (.A(_03900_),
    .B(_03896_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _20222_ (.A(_03898_),
    .B(\core.cpuregs[3][20] ),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2_1 _20223_ (.A(_03901_),
    .B(_03902_),
    .Y(_01267_));
 sky130_fd_sc_hd__buf_6 _20224_ (.A(_09466_),
    .X(_03903_));
 sky130_fd_sc_hd__nand2_1 _20225_ (.A(_03903_),
    .B(_03896_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand2_1 _20226_ (.A(_03898_),
    .B(net180),
    .Y(_03905_));
 sky130_fd_sc_hd__nand2_1 _20227_ (.A(_03904_),
    .B(_03905_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_1 _20228_ (.A(_03720_),
    .B(_03896_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand2_1 _20229_ (.A(_03898_),
    .B(\core.cpuregs[3][22] ),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _20230_ (.A(_03906_),
    .B(_03907_),
    .Y(_01269_));
 sky130_fd_sc_hd__buf_6 _20231_ (.A(_09480_),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_1 _20232_ (.A(_03908_),
    .B(_03896_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand2_1 _20233_ (.A(_03898_),
    .B(\core.cpuregs[3][23] ),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _20234_ (.A(_03909_),
    .B(_03910_),
    .Y(_01270_));
 sky130_fd_sc_hd__buf_6 _20235_ (.A(_09488_),
    .X(_03911_));
 sky130_fd_sc_hd__nand2_1 _20236_ (.A(_03911_),
    .B(_03896_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand2_4 _20237_ (.A(_03898_),
    .B(\core.cpuregs[3][24] ),
    .Y(_03913_));
 sky130_fd_sc_hd__nand2_1 _20238_ (.A(_03912_),
    .B(_03913_),
    .Y(_01271_));
 sky130_fd_sc_hd__clkbuf_2 _20239_ (.A(_09498_),
    .X(_03914_));
 sky130_fd_sc_hd__buf_4 _20240_ (.A(_03856_),
    .X(_03915_));
 sky130_fd_sc_hd__nand2_1 _20241_ (.A(_03914_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20242_ (.A(_03881_),
    .X(_03917_));
 sky130_fd_sc_hd__nand2_1 _20243_ (.A(_03917_),
    .B(\core.cpuregs[3][25] ),
    .Y(_03918_));
 sky130_fd_sc_hd__nand2_1 _20244_ (.A(_03916_),
    .B(_03918_),
    .Y(_01272_));
 sky130_fd_sc_hd__buf_2 _20245_ (.A(_09508_),
    .X(_03919_));
 sky130_fd_sc_hd__nand2_1 _20246_ (.A(_03919_),
    .B(_03915_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand2_1 _20247_ (.A(_03917_),
    .B(\core.cpuregs[3][26] ),
    .Y(_03921_));
 sky130_fd_sc_hd__nand2_1 _20248_ (.A(_03920_),
    .B(_03921_),
    .Y(_01273_));
 sky130_fd_sc_hd__buf_6 _20249_ (.A(_09515_),
    .X(_03922_));
 sky130_fd_sc_hd__nand2_2 _20250_ (.A(_03922_),
    .B(_03915_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_1 _20251_ (.A(_03917_),
    .B(\core.cpuregs[3][27] ),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _20252_ (.A(_03923_),
    .B(_03924_),
    .Y(_01274_));
 sky130_fd_sc_hd__buf_6 _20253_ (.A(_09524_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_1 _20254_ (.A(_03925_),
    .B(_03915_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_1 _20255_ (.A(_03917_),
    .B(net125),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _20256_ (.A(_03926_),
    .B(_03927_),
    .Y(_01275_));
 sky130_fd_sc_hd__buf_4 _20257_ (.A(_09533_),
    .X(_03928_));
 sky130_fd_sc_hd__nand2_4 _20258_ (.A(_03928_),
    .B(_03915_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_2 _20259_ (.A(_03917_),
    .B(\core.cpuregs[3][29] ),
    .Y(_03930_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_03929_),
    .B(_03930_),
    .Y(_01276_));
 sky130_fd_sc_hd__buf_6 _20261_ (.A(_09541_),
    .X(_03931_));
 sky130_fd_sc_hd__nand2_1 _20262_ (.A(_03931_),
    .B(_03915_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _20263_ (.A(_03917_),
    .B(\core.cpuregs[3][30] ),
    .Y(_03933_));
 sky130_fd_sc_hd__nand2_1 _20264_ (.A(_03932_),
    .B(_03933_),
    .Y(_01277_));
 sky130_fd_sc_hd__buf_4 _20265_ (.A(_09550_),
    .X(_03934_));
 sky130_fd_sc_hd__nand2_1 _20266_ (.A(_03934_),
    .B(_03856_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2_1 _20267_ (.A(_03881_),
    .B(\core.cpuregs[3][31] ),
    .Y(_03936_));
 sky130_fd_sc_hd__nand2_1 _20268_ (.A(_03935_),
    .B(_03936_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _20269_ (.A(_03031_),
    .B(_09812_),
    .Y(_03937_));
 sky130_fd_sc_hd__clkbuf_2 _20270_ (.A(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__clkbuf_2 _20271_ (.A(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__mux2_1 _20272_ (.A0(\core.cpuregs[19][0] ),
    .A1(_03853_),
    .S(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__buf_1 _20273_ (.A(_03940_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _20274_ (.A0(\core.cpuregs[19][1] ),
    .A1(_03858_),
    .S(_03939_),
    .X(_03941_));
 sky130_fd_sc_hd__clkbuf_1 _20275_ (.A(_03941_),
    .X(_01280_));
 sky130_fd_sc_hd__clkbuf_4 _20276_ (.A(_03938_),
    .X(_03942_));
 sky130_fd_sc_hd__mux2_1 _20277_ (.A0(\core.cpuregs[19][2] ),
    .A1(_03860_),
    .S(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_1 _20278_ (.A(_03943_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _20279_ (.A0(\core.cpuregs[19][3] ),
    .A1(_03863_),
    .S(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__buf_1 _20280_ (.A(_03944_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _20281_ (.A0(\core.cpuregs[19][4] ),
    .A1(_03865_),
    .S(_03942_),
    .X(_03945_));
 sky130_fd_sc_hd__buf_1 _20282_ (.A(_03945_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _20283_ (.A0(\core.cpuregs[19][5] ),
    .A1(_03867_),
    .S(_03942_),
    .X(_03946_));
 sky130_fd_sc_hd__clkbuf_1 _20284_ (.A(_03946_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _20285_ (.A0(\core.cpuregs[19][6] ),
    .A1(_03869_),
    .S(_03942_),
    .X(_03947_));
 sky130_fd_sc_hd__clkbuf_1 _20286_ (.A(_03947_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _20287_ (.A0(\core.cpuregs[19][7] ),
    .A1(_03871_),
    .S(_03942_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_1 _20288_ (.A(_03948_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _20289_ (.A0(\core.cpuregs[19][8] ),
    .A1(_03873_),
    .S(_03938_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_1 _20290_ (.A(_03949_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _20291_ (.A0(\core.cpuregs[19][9] ),
    .A1(_03875_),
    .S(_03938_),
    .X(_03950_));
 sky130_fd_sc_hd__clkbuf_2 _20292_ (.A(_03950_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _20293_ (.A0(\core.cpuregs[19][10] ),
    .A1(_03877_),
    .S(_03938_),
    .X(_03951_));
 sky130_fd_sc_hd__buf_1 _20294_ (.A(_03951_),
    .X(_01289_));
 sky130_fd_sc_hd__inv_2 _20295_ (.A(_03937_),
    .Y(_03952_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20296_ (.A(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_2 _20297_ (.A0(_03879_),
    .A1(\core.cpuregs[19][11] ),
    .S(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__buf_1 _20298_ (.A(_03954_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _20299_ (.A0(\core.cpuregs[19][12] ),
    .A1(_03883_),
    .S(_03938_),
    .X(_03955_));
 sky130_fd_sc_hd__clkbuf_1 _20300_ (.A(_03955_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _20301_ (.A0(_03885_),
    .A1(\core.cpuregs[19][13] ),
    .S(_03953_),
    .X(_03956_));
 sky130_fd_sc_hd__buf_1 _20302_ (.A(_03956_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _20303_ (.A0(_03887_),
    .A1(\core.cpuregs[19][14] ),
    .S(_03952_),
    .X(_03957_));
 sky130_fd_sc_hd__clkbuf_1 _20304_ (.A(_03957_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _20305_ (.A0(_03889_),
    .A1(\core.cpuregs[19][15] ),
    .S(_03952_),
    .X(_03958_));
 sky130_fd_sc_hd__buf_1 _20306_ (.A(_03958_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_4 _20307_ (.A0(_03891_),
    .A1(\core.cpuregs[19][16] ),
    .S(_03952_),
    .X(_03959_));
 sky130_fd_sc_hd__buf_1 _20308_ (.A(_03959_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _20309_ (.A0(_03893_),
    .A1(\core.cpuregs[19][17] ),
    .S(_03952_),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_1 _20310_ (.A(_03960_),
    .X(_01296_));
 sky130_fd_sc_hd__and2_1 _20311_ (.A(_03953_),
    .B(\core.cpuregs[19][18] ),
    .X(_03961_));
 sky130_fd_sc_hd__a21o_1 _20312_ (.A1(_09442_),
    .A2(_03939_),
    .B1(_03961_),
    .X(_01297_));
 sky130_fd_sc_hd__clkbuf_4 _20313_ (.A(_03939_),
    .X(_03962_));
 sky130_fd_sc_hd__nand2_1 _20314_ (.A(_03711_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20315_ (.A(_03953_),
    .X(_03964_));
 sky130_fd_sc_hd__nand2_2 _20316_ (.A(_03964_),
    .B(\core.cpuregs[19][19] ),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _20317_ (.A(_03963_),
    .B(_03965_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _20318_ (.A(_03900_),
    .B(_03962_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_1 _20319_ (.A(_03964_),
    .B(\core.cpuregs[19][20] ),
    .Y(_03967_));
 sky130_fd_sc_hd__nand2_1 _20320_ (.A(_03966_),
    .B(_03967_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _20321_ (.A(_03903_),
    .B(_03962_),
    .Y(_03968_));
 sky130_fd_sc_hd__nand2_1 _20322_ (.A(_03964_),
    .B(\core.cpuregs[19][21] ),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _20323_ (.A(_03968_),
    .B(_03969_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _20324_ (.A(_03720_),
    .B(_03962_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_03964_),
    .B(\core.cpuregs[19][22] ),
    .Y(_03971_));
 sky130_fd_sc_hd__nand2_1 _20326_ (.A(_03970_),
    .B(_03971_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_2 _20327_ (.A(_03908_),
    .B(_03962_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _20328_ (.A(_03964_),
    .B(\core.cpuregs[19][23] ),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _20329_ (.A(_03972_),
    .B(_03973_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_2 _20330_ (.A(_03911_),
    .B(_03962_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _20331_ (.A(_03964_),
    .B(\core.cpuregs[19][24] ),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _20332_ (.A(_03974_),
    .B(_03975_),
    .Y(_01303_));
 sky130_fd_sc_hd__buf_2 _20333_ (.A(_03939_),
    .X(_03976_));
 sky130_fd_sc_hd__nand2_1 _20334_ (.A(_03914_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__clkbuf_2 _20335_ (.A(_03953_),
    .X(_03978_));
 sky130_fd_sc_hd__nand2_1 _20336_ (.A(_03978_),
    .B(\core.cpuregs[19][25] ),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _20337_ (.A(_03977_),
    .B(_03979_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _20338_ (.A(_03919_),
    .B(_03976_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _20339_ (.A(_03978_),
    .B(\core.cpuregs[19][26] ),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _20340_ (.A(_03980_),
    .B(_03981_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _20341_ (.A(_03922_),
    .B(_03976_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_2 _20342_ (.A(_03978_),
    .B(\core.cpuregs[19][27] ),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _20343_ (.A(_03982_),
    .B(_03983_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_4 _20344_ (.A(_03925_),
    .B(_03976_),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_2 _20345_ (.A(_03978_),
    .B(\core.cpuregs[19][28] ),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _20346_ (.A(_03984_),
    .B(_03985_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _20347_ (.A(_03928_),
    .B(_03976_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _20348_ (.A(_03978_),
    .B(\core.cpuregs[19][29] ),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _20349_ (.A(_03986_),
    .B(_03987_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_4 _20350_ (.A(_03931_),
    .B(_03976_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_1 _20351_ (.A(_03978_),
    .B(\core.cpuregs[19][30] ),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _20352_ (.A(_03988_),
    .B(_03989_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _20353_ (.A(_03934_),
    .B(_03939_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _20354_ (.A(_03953_),
    .B(\core.cpuregs[19][31] ),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _20355_ (.A(_03990_),
    .B(_03991_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _20356_ (.A(_09948_),
    .B(_09812_),
    .Y(_03992_));
 sky130_fd_sc_hd__clkbuf_2 _20357_ (.A(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__clkbuf_2 _20358_ (.A(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _20359_ (.A0(\core.cpuregs[31][0] ),
    .A1(_03853_),
    .S(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20360_ (.A(_03995_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_4 _20361_ (.A0(\core.cpuregs[31][1] ),
    .A1(_03858_),
    .S(_03994_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_1 _20362_ (.A(_03996_),
    .X(_01312_));
 sky130_fd_sc_hd__clkbuf_4 _20363_ (.A(_03993_),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_1 _20364_ (.A0(\core.cpuregs[31][2] ),
    .A1(_03860_),
    .S(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__buf_1 _20365_ (.A(_03998_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _20366_ (.A0(\core.cpuregs[31][3] ),
    .A1(_03863_),
    .S(_03997_),
    .X(_03999_));
 sky130_fd_sc_hd__buf_1 _20367_ (.A(_03999_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _20368_ (.A0(\core.cpuregs[31][4] ),
    .A1(_03865_),
    .S(_03997_),
    .X(_04000_));
 sky130_fd_sc_hd__buf_1 _20369_ (.A(_04000_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _20370_ (.A0(\core.cpuregs[31][5] ),
    .A1(_03867_),
    .S(_03997_),
    .X(_04001_));
 sky130_fd_sc_hd__clkbuf_1 _20371_ (.A(_04001_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _20372_ (.A0(\core.cpuregs[31][6] ),
    .A1(_03869_),
    .S(_03997_),
    .X(_04002_));
 sky130_fd_sc_hd__buf_1 _20373_ (.A(_04002_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_2 _20374_ (.A0(\core.cpuregs[31][7] ),
    .A1(_03871_),
    .S(_03997_),
    .X(_04003_));
 sky130_fd_sc_hd__buf_1 _20375_ (.A(_04003_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _20376_ (.A0(\core.cpuregs[31][8] ),
    .A1(_03873_),
    .S(_03993_),
    .X(_04004_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20377_ (.A(_04004_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _20378_ (.A0(\core.cpuregs[31][9] ),
    .A1(_03875_),
    .S(_03993_),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _20379_ (.A(_04005_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _20380_ (.A0(\core.cpuregs[31][10] ),
    .A1(_03877_),
    .S(_03993_),
    .X(_04006_));
 sky130_fd_sc_hd__buf_1 _20381_ (.A(_04006_),
    .X(_01321_));
 sky130_fd_sc_hd__inv_2 _20382_ (.A(_03992_),
    .Y(_04007_));
 sky130_fd_sc_hd__clkbuf_2 _20383_ (.A(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _20384_ (.A0(_03879_),
    .A1(\core.cpuregs[31][11] ),
    .S(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__buf_1 _20385_ (.A(_04009_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_4 _20386_ (.A0(\core.cpuregs[31][12] ),
    .A1(_03883_),
    .S(_03993_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_1 _20387_ (.A(_04010_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _20388_ (.A0(_03885_),
    .A1(\core.cpuregs[31][13] ),
    .S(_04008_),
    .X(_04011_));
 sky130_fd_sc_hd__buf_1 _20389_ (.A(_04011_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_4 _20390_ (.A0(_03887_),
    .A1(\core.cpuregs[31][14] ),
    .S(_04007_),
    .X(_04012_));
 sky130_fd_sc_hd__clkbuf_1 _20391_ (.A(_04012_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _20392_ (.A0(_03889_),
    .A1(\core.cpuregs[31][15] ),
    .S(_04007_),
    .X(_04013_));
 sky130_fd_sc_hd__clkbuf_1 _20393_ (.A(_04013_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_4 _20394_ (.A0(_03891_),
    .A1(\core.cpuregs[31][16] ),
    .S(_04007_),
    .X(_04014_));
 sky130_fd_sc_hd__buf_1 _20395_ (.A(_04014_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _20396_ (.A0(_03893_),
    .A1(\core.cpuregs[31][17] ),
    .S(_04007_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_1 _20397_ (.A(_04015_),
    .X(_01328_));
 sky130_fd_sc_hd__nand2_1 _20398_ (.A(_04008_),
    .B(\core.cpuregs[31][18] ),
    .Y(_04016_));
 sky130_fd_sc_hd__a21bo_1 _20399_ (.A1(_03198_),
    .A2(_03994_),
    .B1_N(_04016_),
    .X(_01329_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20400_ (.A(_03994_),
    .X(_04017_));
 sky130_fd_sc_hd__nand2_1 _20401_ (.A(_03711_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__clkbuf_4 _20402_ (.A(_04008_),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _20403_ (.A(_04019_),
    .B(net147),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_1 _20404_ (.A(_04018_),
    .B(_04020_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _20405_ (.A(_03900_),
    .B(_04017_),
    .Y(_04021_));
 sky130_fd_sc_hd__nand2_1 _20406_ (.A(_04019_),
    .B(\core.cpuregs[31][20] ),
    .Y(_04022_));
 sky130_fd_sc_hd__nand2_1 _20407_ (.A(_04021_),
    .B(_04022_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _20408_ (.A(_03903_),
    .B(_04017_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(_04019_),
    .B(\core.cpuregs[31][21] ),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _20410_ (.A(_04023_),
    .B(_04024_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _20411_ (.A(_03720_),
    .B(_04017_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _20412_ (.A(_04019_),
    .B(\core.cpuregs[31][22] ),
    .Y(_04026_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(_04025_),
    .B(_04026_),
    .Y(_01333_));
 sky130_fd_sc_hd__nand2_1 _20414_ (.A(_03908_),
    .B(_04017_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand2_1 _20415_ (.A(_04019_),
    .B(\core.cpuregs[31][23] ),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(_04027_),
    .B(_04028_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_2 _20417_ (.A(_03911_),
    .B(_04017_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _20418_ (.A(_04019_),
    .B(\core.cpuregs[31][24] ),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _20419_ (.A(_04029_),
    .B(_04030_),
    .Y(_01335_));
 sky130_fd_sc_hd__clkbuf_4 _20420_ (.A(_03994_),
    .X(_04031_));
 sky130_fd_sc_hd__nand2_1 _20421_ (.A(_03914_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20422_ (.A(_04008_),
    .X(_04033_));
 sky130_fd_sc_hd__nand2_1 _20423_ (.A(_04033_),
    .B(\core.cpuregs[31][25] ),
    .Y(_04034_));
 sky130_fd_sc_hd__nand2_1 _20424_ (.A(_04032_),
    .B(_04034_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _20425_ (.A(_03919_),
    .B(_04031_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _20426_ (.A(_04033_),
    .B(\core.cpuregs[31][26] ),
    .Y(_04036_));
 sky130_fd_sc_hd__nand2_1 _20427_ (.A(_04035_),
    .B(_04036_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _20428_ (.A(_03922_),
    .B(_04031_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2_1 _20429_ (.A(_04033_),
    .B(\core.cpuregs[31][27] ),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_1 _20430_ (.A(_04037_),
    .B(_04038_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _20431_ (.A(_03925_),
    .B(_04031_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_2 _20432_ (.A(_04033_),
    .B(\core.cpuregs[31][28] ),
    .Y(_04040_));
 sky130_fd_sc_hd__nand2_1 _20433_ (.A(_04039_),
    .B(_04040_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2_1 _20434_ (.A(_03928_),
    .B(_04031_),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_1 _20435_ (.A(_04033_),
    .B(\core.cpuregs[31][29] ),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _20436_ (.A(_04041_),
    .B(_04042_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _20437_ (.A(_03931_),
    .B(_04031_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _20438_ (.A(_04033_),
    .B(\core.cpuregs[31][30] ),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _20439_ (.A(_04043_),
    .B(_04044_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_2 _20440_ (.A(_03934_),
    .B(_03994_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_2 _20441_ (.A(_04008_),
    .B(\core.cpuregs[31][31] ),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _20442_ (.A(_04045_),
    .B(_04046_),
    .Y(_01342_));
 sky130_fd_sc_hd__and3_4 _20443_ (.A(_09323_),
    .B(_09557_),
    .C(_10064_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_2 _20444_ (.A(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_2 _20445_ (.A(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__mux2_2 _20446_ (.A0(\core.cpuregs[29][0] ),
    .A1(_03853_),
    .S(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__buf_1 _20447_ (.A(_04050_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _20448_ (.A0(\core.cpuregs[29][1] ),
    .A1(_03858_),
    .S(_04049_),
    .X(_04051_));
 sky130_fd_sc_hd__clkbuf_1 _20449_ (.A(_04051_),
    .X(_01376_));
 sky130_fd_sc_hd__clkbuf_2 _20450_ (.A(_04048_),
    .X(_04052_));
 sky130_fd_sc_hd__mux2_1 _20451_ (.A0(\core.cpuregs[29][2] ),
    .A1(_03860_),
    .S(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__buf_1 _20452_ (.A(_04053_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _20453_ (.A0(\core.cpuregs[29][3] ),
    .A1(_03863_),
    .S(_04052_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_1 _20454_ (.A(_04054_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_2 _20455_ (.A0(\core.cpuregs[29][4] ),
    .A1(_03865_),
    .S(_04052_),
    .X(_04055_));
 sky130_fd_sc_hd__buf_1 _20456_ (.A(_04055_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_2 _20457_ (.A0(\core.cpuregs[29][5] ),
    .A1(_03867_),
    .S(_04052_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _20458_ (.A(_04056_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_2 _20459_ (.A0(\core.cpuregs[29][6] ),
    .A1(_03869_),
    .S(_04052_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _20460_ (.A(_04057_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _20461_ (.A0(\core.cpuregs[29][7] ),
    .A1(_03871_),
    .S(_04052_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _20462_ (.A(_04058_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _20463_ (.A0(\core.cpuregs[29][8] ),
    .A1(_03873_),
    .S(_04048_),
    .X(_04059_));
 sky130_fd_sc_hd__buf_1 _20464_ (.A(_04059_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _20465_ (.A0(\core.cpuregs[29][9] ),
    .A1(_03875_),
    .S(_04048_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _20466_ (.A(_04060_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _20467_ (.A0(\core.cpuregs[29][10] ),
    .A1(_03877_),
    .S(_04048_),
    .X(_04061_));
 sky130_fd_sc_hd__buf_1 _20468_ (.A(_04061_),
    .X(_01385_));
 sky130_fd_sc_hd__inv_2 _20469_ (.A(_04047_),
    .Y(_04062_));
 sky130_fd_sc_hd__buf_2 _20470_ (.A(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__mux2_2 _20471_ (.A0(_03879_),
    .A1(\core.cpuregs[29][11] ),
    .S(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__buf_1 _20472_ (.A(_04064_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _20473_ (.A0(\core.cpuregs[29][12] ),
    .A1(_03883_),
    .S(_04048_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _20474_ (.A(_04065_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _20475_ (.A0(_03885_),
    .A1(\core.cpuregs[29][13] ),
    .S(_04063_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _20476_ (.A(_04066_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _20477_ (.A0(_03887_),
    .A1(\core.cpuregs[29][14] ),
    .S(_04062_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _20478_ (.A(_04067_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _20479_ (.A0(_03889_),
    .A1(\core.cpuregs[29][15] ),
    .S(_04062_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _20480_ (.A(_04068_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _20481_ (.A0(_03891_),
    .A1(\core.cpuregs[29][16] ),
    .S(_04062_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _20482_ (.A(_04069_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _20483_ (.A0(_03893_),
    .A1(\core.cpuregs[29][17] ),
    .S(_04062_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _20484_ (.A(_04070_),
    .X(_01392_));
 sky130_fd_sc_hd__nand2_8 _20485_ (.A(_04063_),
    .B(\core.cpuregs[29][18] ),
    .Y(_04071_));
 sky130_fd_sc_hd__a21bo_1 _20486_ (.A1(_03198_),
    .A2(_04049_),
    .B1_N(_04071_),
    .X(_01393_));
 sky130_fd_sc_hd__clkbuf_2 _20487_ (.A(_04049_),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _20488_ (.A(_03424_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20489_ (.A(_04063_),
    .X(_04074_));
 sky130_fd_sc_hd__nand2_1 _20490_ (.A(_04074_),
    .B(\core.cpuregs[29][19] ),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _20491_ (.A(_04073_),
    .B(_04075_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_4 _20492_ (.A(_03900_),
    .B(_04072_),
    .Y(_04076_));
 sky130_fd_sc_hd__nand2_2 _20493_ (.A(_04074_),
    .B(\core.cpuregs[29][20] ),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _20494_ (.A(_04076_),
    .B(_04077_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _20495_ (.A(_03903_),
    .B(_04072_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _20496_ (.A(_04074_),
    .B(net138),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _20497_ (.A(_04078_),
    .B(_04079_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _20498_ (.A(_03435_),
    .B(_04072_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _20499_ (.A(_04074_),
    .B(\core.cpuregs[29][22] ),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_1 _20500_ (.A(_04080_),
    .B(_04081_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _20501_ (.A(_03908_),
    .B(_04072_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _20502_ (.A(_04074_),
    .B(\core.cpuregs[29][23] ),
    .Y(_04083_));
 sky130_fd_sc_hd__nand2_1 _20503_ (.A(_04082_),
    .B(_04083_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _20504_ (.A(_03911_),
    .B(_04072_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _20505_ (.A(_04074_),
    .B(\core.cpuregs[29][24] ),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _20506_ (.A(_04084_),
    .B(_04085_),
    .Y(_01399_));
 sky130_fd_sc_hd__clkbuf_4 _20507_ (.A(_04049_),
    .X(_04086_));
 sky130_fd_sc_hd__nand2_1 _20508_ (.A(_03914_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20509_ (.A(_04063_),
    .X(_04088_));
 sky130_fd_sc_hd__nand2_1 _20510_ (.A(_04088_),
    .B(\core.cpuregs[29][25] ),
    .Y(_04089_));
 sky130_fd_sc_hd__nand2_1 _20511_ (.A(_04087_),
    .B(_04089_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_1 _20512_ (.A(_03919_),
    .B(_04086_),
    .Y(_04090_));
 sky130_fd_sc_hd__nand2_1 _20513_ (.A(_04088_),
    .B(\core.cpuregs[29][26] ),
    .Y(_04091_));
 sky130_fd_sc_hd__nand2_1 _20514_ (.A(_04090_),
    .B(_04091_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand2_2 _20515_ (.A(_03922_),
    .B(_04086_),
    .Y(_04092_));
 sky130_fd_sc_hd__nand2_1 _20516_ (.A(_04088_),
    .B(\core.cpuregs[29][27] ),
    .Y(_04093_));
 sky130_fd_sc_hd__nand2_1 _20517_ (.A(_04092_),
    .B(_04093_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_1 _20518_ (.A(_03925_),
    .B(_04086_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _20519_ (.A(_04088_),
    .B(\core.cpuregs[29][28] ),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_1 _20520_ (.A(_04094_),
    .B(_04095_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand2_2 _20521_ (.A(_03928_),
    .B(_04086_),
    .Y(_04096_));
 sky130_fd_sc_hd__nand2_2 _20522_ (.A(_04088_),
    .B(\core.cpuregs[29][29] ),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_1 _20523_ (.A(_04096_),
    .B(_04097_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_2 _20524_ (.A(_03931_),
    .B(_04086_),
    .Y(_04098_));
 sky130_fd_sc_hd__nand2_1 _20525_ (.A(_04088_),
    .B(\core.cpuregs[29][30] ),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _20526_ (.A(_04098_),
    .B(_04099_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand2_1 _20527_ (.A(_03934_),
    .B(_04049_),
    .Y(_04100_));
 sky130_fd_sc_hd__nand2_1 _20528_ (.A(_04063_),
    .B(\core.cpuregs[29][31] ),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _20529_ (.A(_04100_),
    .B(_04101_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _20530_ (.A(_03031_),
    .B(_10158_),
    .Y(_04102_));
 sky130_fd_sc_hd__clkbuf_2 _20531_ (.A(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_2 _20532_ (.A(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__mux2_1 _20533_ (.A0(\core.cpuregs[18][0] ),
    .A1(_03853_),
    .S(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _20534_ (.A(_04105_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _20535_ (.A0(\core.cpuregs[18][1] ),
    .A1(_03858_),
    .S(_04104_),
    .X(_04106_));
 sky130_fd_sc_hd__buf_1 _20536_ (.A(_04106_),
    .X(_01408_));
 sky130_fd_sc_hd__clkbuf_4 _20537_ (.A(_04103_),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _20538_ (.A0(\core.cpuregs[18][2] ),
    .A1(_03860_),
    .S(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__buf_1 _20539_ (.A(_04108_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _20540_ (.A0(\core.cpuregs[18][3] ),
    .A1(_03863_),
    .S(_04107_),
    .X(_04109_));
 sky130_fd_sc_hd__buf_1 _20541_ (.A(_04109_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _20542_ (.A0(\core.cpuregs[18][4] ),
    .A1(_03865_),
    .S(_04107_),
    .X(_04110_));
 sky130_fd_sc_hd__buf_1 _20543_ (.A(_04110_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _20544_ (.A0(\core.cpuregs[18][5] ),
    .A1(_03867_),
    .S(_04107_),
    .X(_04111_));
 sky130_fd_sc_hd__buf_1 _20545_ (.A(_04111_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_2 _20546_ (.A0(\core.cpuregs[18][6] ),
    .A1(_03869_),
    .S(_04107_),
    .X(_04112_));
 sky130_fd_sc_hd__buf_1 _20547_ (.A(_04112_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _20548_ (.A0(\core.cpuregs[18][7] ),
    .A1(_03871_),
    .S(_04107_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _20549_ (.A(_04113_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _20550_ (.A0(\core.cpuregs[18][8] ),
    .A1(_03873_),
    .S(_04103_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _20551_ (.A(_04114_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _20552_ (.A0(\core.cpuregs[18][9] ),
    .A1(_03875_),
    .S(_04103_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _20553_ (.A(_04115_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _20554_ (.A0(\core.cpuregs[18][10] ),
    .A1(_03877_),
    .S(_04103_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _20555_ (.A(_04116_),
    .X(_01417_));
 sky130_fd_sc_hd__inv_2 _20556_ (.A(_04102_),
    .Y(_04117_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20557_ (.A(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__mux2_1 _20558_ (.A0(_03879_),
    .A1(\core.cpuregs[18][11] ),
    .S(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _20559_ (.A(_04119_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_8 _20560_ (.A0(\core.cpuregs[18][12] ),
    .A1(_03883_),
    .S(_04103_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _20561_ (.A(_04120_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _20562_ (.A0(_03885_),
    .A1(\core.cpuregs[18][13] ),
    .S(_04118_),
    .X(_04121_));
 sky130_fd_sc_hd__buf_1 _20563_ (.A(_04121_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_4 _20564_ (.A0(_03887_),
    .A1(\core.cpuregs[18][14] ),
    .S(_04117_),
    .X(_04122_));
 sky130_fd_sc_hd__buf_1 _20565_ (.A(_04122_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _20566_ (.A0(_03889_),
    .A1(\core.cpuregs[18][15] ),
    .S(_04117_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _20567_ (.A(_04123_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _20568_ (.A0(_03891_),
    .A1(\core.cpuregs[18][16] ),
    .S(_04117_),
    .X(_04124_));
 sky130_fd_sc_hd__buf_4 _20569_ (.A(_04124_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _20570_ (.A0(_03893_),
    .A1(\core.cpuregs[18][17] ),
    .S(_04117_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _20571_ (.A(_04125_),
    .X(_01424_));
 sky130_fd_sc_hd__and2_1 _20572_ (.A(_04118_),
    .B(\core.cpuregs[18][18] ),
    .X(_04126_));
 sky130_fd_sc_hd__a21o_1 _20573_ (.A1(_09442_),
    .A2(_04104_),
    .B1(_04126_),
    .X(_01425_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20574_ (.A(_04104_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_1 _20575_ (.A(_03424_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__clkbuf_4 _20576_ (.A(_04118_),
    .X(_04129_));
 sky130_fd_sc_hd__nand2_1 _20577_ (.A(_04129_),
    .B(\core.cpuregs[18][19] ),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _20578_ (.A(_04128_),
    .B(_04130_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _20579_ (.A(_03900_),
    .B(_04127_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _20580_ (.A(_04129_),
    .B(\core.cpuregs[18][20] ),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _20581_ (.A(_04131_),
    .B(_04132_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _20582_ (.A(_03903_),
    .B(_04127_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand2_1 _20583_ (.A(_04129_),
    .B(net164),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _20584_ (.A(_04133_),
    .B(_04134_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _20585_ (.A(_03435_),
    .B(_04127_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand2_1 _20586_ (.A(_04129_),
    .B(\core.cpuregs[18][22] ),
    .Y(_04136_));
 sky130_fd_sc_hd__nand2_1 _20587_ (.A(_04135_),
    .B(_04136_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _20588_ (.A(_03908_),
    .B(_04127_),
    .Y(_04137_));
 sky130_fd_sc_hd__nand2_1 _20589_ (.A(_04129_),
    .B(\core.cpuregs[18][23] ),
    .Y(_04138_));
 sky130_fd_sc_hd__nand2_1 _20590_ (.A(_04137_),
    .B(_04138_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _20591_ (.A(_03911_),
    .B(_04127_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _20592_ (.A(_04129_),
    .B(net121),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2_1 _20593_ (.A(_04139_),
    .B(_04140_),
    .Y(_01431_));
 sky130_fd_sc_hd__clkbuf_4 _20594_ (.A(_04104_),
    .X(_04141_));
 sky130_fd_sc_hd__nand2_1 _20595_ (.A(_03914_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__clkbuf_2 _20596_ (.A(_04118_),
    .X(_04143_));
 sky130_fd_sc_hd__nand2_1 _20597_ (.A(_04143_),
    .B(\core.cpuregs[18][25] ),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _20598_ (.A(_04142_),
    .B(_04144_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _20599_ (.A(_03919_),
    .B(_04141_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _20600_ (.A(_04143_),
    .B(\core.cpuregs[18][26] ),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_1 _20601_ (.A(_04145_),
    .B(_04146_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _20602_ (.A(_03922_),
    .B(_04141_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _20603_ (.A(_04143_),
    .B(net184),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _20604_ (.A(_04147_),
    .B(_04148_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _20605_ (.A(_03925_),
    .B(_04141_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_1 _20606_ (.A(_04143_),
    .B(\core.cpuregs[18][28] ),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _20607_ (.A(_04149_),
    .B(_04150_),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _20608_ (.A(_03928_),
    .B(_04141_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_1 _20609_ (.A(_04143_),
    .B(\core.cpuregs[18][29] ),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2_1 _20610_ (.A(_04151_),
    .B(_04152_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _20611_ (.A(_03931_),
    .B(_04141_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand2_4 _20612_ (.A(_04143_),
    .B(\core.cpuregs[18][30] ),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _20613_ (.A(_04153_),
    .B(_04154_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _20614_ (.A(_03934_),
    .B(_04104_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _20615_ (.A(_04118_),
    .B(\core.cpuregs[18][31] ),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _20616_ (.A(_04155_),
    .B(_04156_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _20617_ (.A(_09811_),
    .B(_09949_),
    .Y(_04157_));
 sky130_fd_sc_hd__buf_4 _20618_ (.A(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_2 _20619_ (.A(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__mux2_1 _20620_ (.A0(\core.cpuregs[24][0] ),
    .A1(_03853_),
    .S(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__buf_1 _20621_ (.A(_04160_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_4 _20622_ (.A0(\core.cpuregs[24][1] ),
    .A1(_03858_),
    .S(_04159_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _20623_ (.A(_04161_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_4 _20624_ (.A(_04158_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _20625_ (.A0(\core.cpuregs[24][2] ),
    .A1(_03860_),
    .S(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__buf_1 _20626_ (.A(_04163_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _20627_ (.A0(\core.cpuregs[24][3] ),
    .A1(_03863_),
    .S(_04162_),
    .X(_04164_));
 sky130_fd_sc_hd__buf_1 _20628_ (.A(_04164_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_4 _20629_ (.A0(\core.cpuregs[24][4] ),
    .A1(_03865_),
    .S(_04162_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _20630_ (.A(_04165_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_2 _20631_ (.A0(\core.cpuregs[24][5] ),
    .A1(_03867_),
    .S(_04162_),
    .X(_04166_));
 sky130_fd_sc_hd__buf_1 _20632_ (.A(_04166_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _20633_ (.A0(\core.cpuregs[24][6] ),
    .A1(_03869_),
    .S(_04162_),
    .X(_04167_));
 sky130_fd_sc_hd__buf_1 _20634_ (.A(_04167_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _20635_ (.A0(\core.cpuregs[24][7] ),
    .A1(_03871_),
    .S(_04162_),
    .X(_04168_));
 sky130_fd_sc_hd__buf_1 _20636_ (.A(_04168_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _20637_ (.A0(\core.cpuregs[24][8] ),
    .A1(_03873_),
    .S(_04158_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _20638_ (.A(_04169_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _20639_ (.A0(\core.cpuregs[24][9] ),
    .A1(_03875_),
    .S(_04158_),
    .X(_04170_));
 sky130_fd_sc_hd__buf_1 _20640_ (.A(_04170_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _20641_ (.A0(\core.cpuregs[24][10] ),
    .A1(_03877_),
    .S(_04158_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _20642_ (.A(_04171_),
    .X(_01449_));
 sky130_fd_sc_hd__inv_2 _20643_ (.A(_04157_),
    .Y(_04172_));
 sky130_fd_sc_hd__clkbuf_2 _20644_ (.A(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__mux2_4 _20645_ (.A0(_03879_),
    .A1(\core.cpuregs[24][11] ),
    .S(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _20646_ (.A(_04174_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_2 _20647_ (.A0(\core.cpuregs[24][12] ),
    .A1(_03883_),
    .S(_04158_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _20648_ (.A(_04175_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _20649_ (.A0(_03885_),
    .A1(\core.cpuregs[24][13] ),
    .S(_04173_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _20650_ (.A(_04176_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_4 _20651_ (.A0(_03887_),
    .A1(\core.cpuregs[24][14] ),
    .S(_04172_),
    .X(_04177_));
 sky130_fd_sc_hd__buf_1 _20652_ (.A(_04177_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _20653_ (.A0(_03889_),
    .A1(\core.cpuregs[24][15] ),
    .S(_04172_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _20654_ (.A(_04178_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _20655_ (.A0(_03891_),
    .A1(\core.cpuregs[24][16] ),
    .S(_04172_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _20656_ (.A(_04179_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _20657_ (.A0(_03893_),
    .A1(\core.cpuregs[24][17] ),
    .S(_04172_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _20658_ (.A(_04180_),
    .X(_01456_));
 sky130_fd_sc_hd__nand2_1 _20659_ (.A(_04173_),
    .B(\core.cpuregs[24][18] ),
    .Y(_04181_));
 sky130_fd_sc_hd__a21bo_1 _20660_ (.A1(_09441_),
    .A2(_04159_),
    .B1_N(_04181_),
    .X(_01457_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20661_ (.A(_04159_),
    .X(_04182_));
 sky130_fd_sc_hd__nand2_1 _20662_ (.A(_03424_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20663_ (.A(_04173_),
    .X(_04184_));
 sky130_fd_sc_hd__nand2_1 _20664_ (.A(_04184_),
    .B(\core.cpuregs[24][19] ),
    .Y(_04185_));
 sky130_fd_sc_hd__nand2_1 _20665_ (.A(_04183_),
    .B(_04185_),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_2 _20666_ (.A(_03900_),
    .B(_04182_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_1 _20667_ (.A(_04184_),
    .B(net181),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_1 _20668_ (.A(_04186_),
    .B(_04187_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_1 _20669_ (.A(_03903_),
    .B(_04182_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _20670_ (.A(_04184_),
    .B(net177),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _20671_ (.A(_04188_),
    .B(_04189_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _20672_ (.A(_03435_),
    .B(_04182_),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _20673_ (.A(_04184_),
    .B(\core.cpuregs[24][22] ),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _20674_ (.A(_04190_),
    .B(_04191_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _20675_ (.A(_03908_),
    .B(_04182_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_1 _20676_ (.A(_04184_),
    .B(\core.cpuregs[24][23] ),
    .Y(_04193_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_04192_),
    .B(_04193_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _20678_ (.A(_03911_),
    .B(_04182_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _20679_ (.A(_04184_),
    .B(\core.cpuregs[24][24] ),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _20680_ (.A(_04194_),
    .B(_04195_),
    .Y(_01463_));
 sky130_fd_sc_hd__clkbuf_2 _20681_ (.A(_04159_),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_4 _20682_ (.A(_03914_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__clkbuf_2 _20683_ (.A(_04173_),
    .X(_04198_));
 sky130_fd_sc_hd__nand2_4 _20684_ (.A(_04198_),
    .B(\core.cpuregs[24][25] ),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _20685_ (.A(_04197_),
    .B(_04199_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _20686_ (.A(_03919_),
    .B(_04196_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _20687_ (.A(_04198_),
    .B(\core.cpuregs[24][26] ),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2_1 _20688_ (.A(_04200_),
    .B(_04201_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _20689_ (.A(_03922_),
    .B(_04196_),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_1 _20690_ (.A(_04198_),
    .B(\core.cpuregs[24][27] ),
    .Y(_04203_));
 sky130_fd_sc_hd__nand2_1 _20691_ (.A(_04202_),
    .B(_04203_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_2 _20692_ (.A(_03925_),
    .B(_04196_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_1 _20693_ (.A(_04198_),
    .B(\core.cpuregs[24][28] ),
    .Y(_04205_));
 sky130_fd_sc_hd__nand2_1 _20694_ (.A(_04204_),
    .B(_04205_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _20695_ (.A(_03928_),
    .B(_04196_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand2_1 _20696_ (.A(_04198_),
    .B(\core.cpuregs[24][29] ),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_4 _20697_ (.A(_04206_),
    .B(_04207_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _20698_ (.A(_03931_),
    .B(_04196_),
    .Y(_04208_));
 sky130_fd_sc_hd__nand2_2 _20699_ (.A(_04198_),
    .B(\core.cpuregs[24][30] ),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _20700_ (.A(_04208_),
    .B(_04209_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_4 _20701_ (.A(_03934_),
    .B(_04159_),
    .Y(_04210_));
 sky130_fd_sc_hd__nand2_1 _20702_ (.A(_04173_),
    .B(net169),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_1 _20703_ (.A(_04210_),
    .B(_04211_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _20704_ (.A(_03396_),
    .B(_02778_),
    .Y(_04212_));
 sky130_fd_sc_hd__clkbuf_4 _20705_ (.A(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_2 _20706_ (.A(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_2 _20707_ (.A0(\core.cpuregs[9][0] ),
    .A1(_09314_),
    .S(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _20708_ (.A(_04215_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _20709_ (.A0(\core.cpuregs[9][1] ),
    .A1(_09336_),
    .S(_04214_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_4 _20710_ (.A(_04216_),
    .X(_01472_));
 sky130_fd_sc_hd__clkbuf_4 _20711_ (.A(_04213_),
    .X(_04217_));
 sky130_fd_sc_hd__mux2_1 _20712_ (.A0(\core.cpuregs[9][2] ),
    .A1(_09339_),
    .S(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__buf_1 _20713_ (.A(_04218_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _20714_ (.A0(\core.cpuregs[9][3] ),
    .A1(_09348_),
    .S(_04217_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _20715_ (.A(_04219_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _20716_ (.A0(\core.cpuregs[9][4] ),
    .A1(_09356_),
    .S(_04217_),
    .X(_04220_));
 sky130_fd_sc_hd__buf_1 _20717_ (.A(_04220_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _20718_ (.A0(\core.cpuregs[9][5] ),
    .A1(_09362_),
    .S(_04217_),
    .X(_04221_));
 sky130_fd_sc_hd__buf_1 _20719_ (.A(_04221_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _20720_ (.A0(\core.cpuregs[9][6] ),
    .A1(_09368_),
    .S(_04217_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _20721_ (.A(_04222_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _20722_ (.A0(\core.cpuregs[9][7] ),
    .A1(_09374_),
    .S(_04217_),
    .X(_04223_));
 sky130_fd_sc_hd__buf_1 _20723_ (.A(_04223_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _20724_ (.A0(\core.cpuregs[9][8] ),
    .A1(_09380_),
    .S(_04213_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _20725_ (.A(_04224_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _20726_ (.A0(\core.cpuregs[9][9] ),
    .A1(_09387_),
    .S(_04213_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _20727_ (.A(_04225_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _20728_ (.A0(\core.cpuregs[9][10] ),
    .A1(_09394_),
    .S(_04213_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _20729_ (.A(_04226_),
    .X(_01481_));
 sky130_fd_sc_hd__inv_2 _20730_ (.A(_04212_),
    .Y(_04227_));
 sky130_fd_sc_hd__clkbuf_2 _20731_ (.A(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__mux2_8 _20732_ (.A0(_09400_),
    .A1(\core.cpuregs[9][11] ),
    .S(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_2 _20733_ (.A(_04229_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _20734_ (.A0(\core.cpuregs[9][12] ),
    .A1(_09407_),
    .S(_04213_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _20735_ (.A(_04230_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _20736_ (.A0(_09413_),
    .A1(\core.cpuregs[9][13] ),
    .S(_04228_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _20737_ (.A(_04231_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_8 _20738_ (.A0(_09418_),
    .A1(\core.cpuregs[9][14] ),
    .S(_04227_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _20739_ (.A(_04232_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _20740_ (.A0(_09423_),
    .A1(\core.cpuregs[9][15] ),
    .S(_04227_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _20741_ (.A(_04233_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _20742_ (.A0(_09430_),
    .A1(\core.cpuregs[9][16] ),
    .S(_04227_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_2 _20743_ (.A(_04234_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _20744_ (.A0(_09435_),
    .A1(\core.cpuregs[9][17] ),
    .S(_04227_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _20745_ (.A(_04235_),
    .X(_01488_));
 sky130_fd_sc_hd__and2_1 _20746_ (.A(_04228_),
    .B(\core.cpuregs[9][18] ),
    .X(_04236_));
 sky130_fd_sc_hd__a21o_1 _20747_ (.A1(_09442_),
    .A2(_04214_),
    .B1(_04236_),
    .X(_01489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20748_ (.A(_04214_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _20749_ (.A(_03424_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__buf_2 _20750_ (.A(_04228_),
    .X(_04239_));
 sky130_fd_sc_hd__nand2_1 _20751_ (.A(_04239_),
    .B(\core.cpuregs[9][19] ),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _20752_ (.A(_04238_),
    .B(_04240_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _20753_ (.A(_09457_),
    .B(_04237_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_1 _20754_ (.A(_04239_),
    .B(\core.cpuregs[9][20] ),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2_1 _20755_ (.A(_04241_),
    .B(_04242_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _20756_ (.A(_09466_),
    .B(_04237_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _20757_ (.A(_04239_),
    .B(net168),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _20758_ (.A(_04243_),
    .B(_04244_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _20759_ (.A(_03435_),
    .B(_04237_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_1 _20760_ (.A(_04239_),
    .B(\core.cpuregs[9][22] ),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _20761_ (.A(_04245_),
    .B(_04246_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _20762_ (.A(_09480_),
    .B(_04237_),
    .Y(_04247_));
 sky130_fd_sc_hd__nand2_1 _20763_ (.A(_04239_),
    .B(net171),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_1 _20764_ (.A(_04247_),
    .B(_04248_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _20765_ (.A(_09488_),
    .B(_04237_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _20766_ (.A(_04239_),
    .B(net154),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _20767_ (.A(_04249_),
    .B(_04250_),
    .Y(_01495_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20768_ (.A(_04214_),
    .X(_04251_));
 sky130_fd_sc_hd__nand2_1 _20769_ (.A(_09498_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _20770_ (.A(_04228_),
    .X(_04253_));
 sky130_fd_sc_hd__nand2_1 _20771_ (.A(_04253_),
    .B(\core.cpuregs[9][25] ),
    .Y(_04254_));
 sky130_fd_sc_hd__nand2_1 _20772_ (.A(_04252_),
    .B(_04254_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _20773_ (.A(_09508_),
    .B(_04251_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_2 _20774_ (.A(_04253_),
    .B(\core.cpuregs[9][26] ),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2_1 _20775_ (.A(_04255_),
    .B(_04256_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(_09515_),
    .B(_04251_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(_04253_),
    .B(\core.cpuregs[9][27] ),
    .Y(_04258_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(_04257_),
    .B(_04258_),
    .Y(_01498_));
 sky130_fd_sc_hd__nand2_1 _20779_ (.A(_09524_),
    .B(_04251_),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _20780_ (.A(_04253_),
    .B(net182),
    .Y(_04260_));
 sky130_fd_sc_hd__nand2_1 _20781_ (.A(_04259_),
    .B(_04260_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _20782_ (.A(_09533_),
    .B(_04251_),
    .Y(_04261_));
 sky130_fd_sc_hd__nand2_1 _20783_ (.A(_04253_),
    .B(net191),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_1 _20784_ (.A(_04261_),
    .B(_04262_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_09541_),
    .B(_04251_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_1 _20786_ (.A(_04253_),
    .B(net150),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_1 _20787_ (.A(_04263_),
    .B(_04264_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand2_1 _20788_ (.A(_09550_),
    .B(_04214_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _20789_ (.A(_04228_),
    .B(\core.cpuregs[9][31] ),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2_1 _20790_ (.A(_04265_),
    .B(_04266_),
    .Y(_01502_));
 sky130_fd_sc_hd__a22o_1 _20791_ (.A1(\core.instr_lhu ),
    .A2(_10218_),
    .B1(_10249_),
    .B2(_02722_),
    .X(_01503_));
 sky130_fd_sc_hd__a22o_1 _20792_ (.A1(\core.instr_lbu ),
    .A2(_10218_),
    .B1(_10260_),
    .B2(_02722_),
    .X(_01504_));
 sky130_fd_sc_hd__a22o_1 _20793_ (.A1(\core.instr_lw ),
    .A2(_10218_),
    .B1(_10222_),
    .B2(_02722_),
    .X(_01505_));
 sky130_fd_sc_hd__a22o_1 _20794_ (.A1(\core.instr_lh ),
    .A2(_10306_),
    .B1(_02722_),
    .B2(_10059_),
    .X(_01506_));
 sky130_fd_sc_hd__or3_2 _20795_ (.A(_10153_),
    .B(_10057_),
    .C(_10154_),
    .X(_04267_));
 sky130_fd_sc_hd__o22a_1 _20796_ (.A1(_04434_),
    .A2(_10054_),
    .B1(_10056_),
    .B2(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__nor2_1 _20797_ (.A(_06372_),
    .B(_04268_),
    .Y(_01507_));
 sky130_fd_sc_hd__o2bb2a_1 _20798_ (.A1_N(\core.instr_blt ),
    .A2_N(_10226_),
    .B1(_10056_),
    .B2(_10261_),
    .X(_04269_));
 sky130_fd_sc_hd__nor2_1 _20799_ (.A(_06372_),
    .B(_04269_),
    .Y(_01508_));
 sky130_fd_sc_hd__or4_2 _20800_ (.A(\core.mem_rdata_q[22] ),
    .B(\core.mem_rdata_q[23] ),
    .C(_10302_),
    .D(\core.mem_rdata_q[20] ),
    .X(_04270_));
 sky130_fd_sc_hd__nor2_1 _20801_ (.A(_10217_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__a32o_1 _20802_ (.A1(_10296_),
    .A2(_10301_),
    .A3(_04271_),
    .B1(_05087_),
    .B2(_10306_),
    .X(_01509_));
 sky130_fd_sc_hd__and2_1 _20803_ (.A(_10292_),
    .B(_10301_),
    .X(_04272_));
 sky130_fd_sc_hd__and3_1 _20804_ (.A(_10239_),
    .B(_10293_),
    .C(_10240_),
    .X(_04273_));
 sky130_fd_sc_hd__a32o_1 _20805_ (.A1(_04272_),
    .A2(_04271_),
    .A3(_04273_),
    .B1(_05042_),
    .B2(_10306_),
    .X(_01510_));
 sky130_fd_sc_hd__a32o_1 _20806_ (.A1(_04272_),
    .A2(_10305_),
    .A3(_04273_),
    .B1(net110),
    .B2(_10254_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_1 _20807_ (.A(_10217_),
    .B(\core.instr_srai ),
    .X(_04274_));
 sky130_fd_sc_hd__a31o_1 _20808_ (.A1(_10268_),
    .A2(_10247_),
    .A3(_10250_),
    .B1(_04274_),
    .X(_01512_));
 sky130_fd_sc_hd__or3_1 _20809_ (.A(_10257_),
    .B(_04267_),
    .C(_10245_),
    .X(_04275_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(_10312_),
    .B(\core.instr_and ),
    .Y(_04276_));
 sky130_fd_sc_hd__buf_2 _20811_ (.A(_04514_),
    .X(_04277_));
 sky130_fd_sc_hd__a21oi_1 _20812_ (.A1(_04275_),
    .A2(_04276_),
    .B1(_04277_),
    .Y(_01513_));
 sky130_fd_sc_hd__or3_1 _20813_ (.A(_10229_),
    .B(_10257_),
    .C(_10244_),
    .X(_04278_));
 sky130_fd_sc_hd__nand2_1 _20814_ (.A(_10312_),
    .B(\core.instr_or ),
    .Y(_04279_));
 sky130_fd_sc_hd__a21oi_1 _20815_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04277_),
    .Y(_01514_));
 sky130_fd_sc_hd__or3_1 _20816_ (.A(_10225_),
    .B(_10264_),
    .C(_10244_),
    .X(_04280_));
 sky130_fd_sc_hd__nand2_1 _20817_ (.A(_10312_),
    .B(\core.instr_srl ),
    .Y(_04281_));
 sky130_fd_sc_hd__a21oi_1 _20818_ (.A1(_04280_),
    .A2(_04281_),
    .B1(_04277_),
    .Y(_01515_));
 sky130_fd_sc_hd__or3_1 _20819_ (.A(_10227_),
    .B(_10257_),
    .C(_10244_),
    .X(_04282_));
 sky130_fd_sc_hd__nand2_1 _20820_ (.A(_10312_),
    .B(\core.instr_sltu ),
    .Y(_04283_));
 sky130_fd_sc_hd__a21oi_1 _20821_ (.A1(_04282_),
    .A2(_04283_),
    .B1(_04277_),
    .Y(_01516_));
 sky130_fd_sc_hd__or3_1 _20822_ (.A(_10223_),
    .B(_10257_),
    .C(_10244_),
    .X(_04284_));
 sky130_fd_sc_hd__nand2_1 _20823_ (.A(_10312_),
    .B(\core.instr_slt ),
    .Y(_04285_));
 sky130_fd_sc_hd__a21oi_1 _20824_ (.A1(_04284_),
    .A2(_04285_),
    .B1(_04277_),
    .Y(_01517_));
 sky130_fd_sc_hd__or3_1 _20825_ (.A(_10225_),
    .B(_10252_),
    .C(_10269_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(_10217_),
    .B(_05802_),
    .Y(_04287_));
 sky130_fd_sc_hd__a21oi_1 _20827_ (.A1(_04286_),
    .A2(_04287_),
    .B1(_04277_),
    .Y(_01518_));
 sky130_fd_sc_hd__a32o_1 _20828_ (.A1(_10246_),
    .A2(_10059_),
    .A3(_02940_),
    .B1(net119),
    .B2(_10254_),
    .X(_01519_));
 sky130_fd_sc_hd__a22o_1 _20829_ (.A1(\core.instr_sw ),
    .A2(_10306_),
    .B1(_10222_),
    .B2(_10220_),
    .X(_01520_));
 sky130_fd_sc_hd__o2bb2a_1 _20830_ (.A1_N(\core.instr_andi ),
    .A2_N(_10216_),
    .B1(_10221_),
    .B2(_04267_),
    .X(_04288_));
 sky130_fd_sc_hd__nor2_1 _20831_ (.A(_06372_),
    .B(_04288_),
    .Y(_01521_));
 sky130_fd_sc_hd__a22o_1 _20832_ (.A1(\core.instr_xori ),
    .A2(_10216_),
    .B1(_10260_),
    .B2(_02940_),
    .X(_04289_));
 sky130_fd_sc_hd__and2_1 _20833_ (.A(_04289_),
    .B(_06506_),
    .X(_04290_));
 sky130_fd_sc_hd__buf_1 _20834_ (.A(_04290_),
    .X(_01522_));
 sky130_fd_sc_hd__a22o_1 _20835_ (.A1(\core.instr_addi ),
    .A2(_10216_),
    .B1(_10155_),
    .B2(_02940_),
    .X(_04291_));
 sky130_fd_sc_hd__and2_1 _20836_ (.A(_04291_),
    .B(_06329_),
    .X(_04292_));
 sky130_fd_sc_hd__buf_1 _20837_ (.A(_04292_),
    .X(_01523_));
 sky130_fd_sc_hd__a22o_1 _20838_ (.A1(\core.instr_sb ),
    .A2(_10306_),
    .B1(_10155_),
    .B2(_10220_),
    .X(_01524_));
 sky130_fd_sc_hd__o21ai_1 _20839_ (.A1(_04369_),
    .A2(_10316_),
    .B1(_04407_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _20840_ (.A(_04472_),
    .B(_04465_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand2_1 _20841_ (.A(_04474_),
    .B(\core.is_sll_srl_sra ),
    .Y(_04294_));
 sky130_fd_sc_hd__nand3_1 _20842_ (.A(_04464_),
    .B(_04466_),
    .C(_10317_),
    .Y(_04295_));
 sky130_fd_sc_hd__nor3_1 _20843_ (.A(_04293_),
    .B(_04294_),
    .C(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__nand2_1 _20844_ (.A(_04293_),
    .B(_04466_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _20845_ (.A(_10317_),
    .B(_10233_),
    .Y(_04298_));
 sky130_fd_sc_hd__o22a_1 _20846_ (.A1(_04484_),
    .A2(_10316_),
    .B1(_04632_),
    .B2(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__o21ai_2 _20847_ (.A1(_10316_),
    .A2(_04297_),
    .B1(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__nor2_1 _20848_ (.A(_04296_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand2_2 _20849_ (.A(_10314_),
    .B(_06316_),
    .Y(_04302_));
 sky130_fd_sc_hd__or2_1 _20850_ (.A(_04302_),
    .B(_04976_),
    .X(_04303_));
 sky130_fd_sc_hd__nand2_1 _20851_ (.A(_04474_),
    .B(_04468_),
    .Y(_04304_));
 sky130_fd_sc_hd__a31o_1 _20852_ (.A1(_04464_),
    .A2(_04367_),
    .A3(_04304_),
    .B1(_04439_),
    .X(_04305_));
 sky130_fd_sc_hd__a21oi_1 _20853_ (.A1(\core.mem_do_prefetch ),
    .A2(_05115_),
    .B1(_06314_),
    .Y(_04306_));
 sky130_fd_sc_hd__o21ai_1 _20854_ (.A1(_04503_),
    .A2(_06315_),
    .B1(_10317_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_1 _20855_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__nand2_1 _20856_ (.A(_04308_),
    .B(_04301_),
    .Y(_04309_));
 sky130_fd_sc_hd__o211ai_2 _20857_ (.A1(_04368_),
    .A2(_04301_),
    .B1(_04303_),
    .C1(_04309_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_4 _20858_ (.A(_04502_),
    .B(_06636_),
    .Y(_04310_));
 sky130_fd_sc_hd__mux2_1 _20859_ (.A0(_04425_),
    .A1(\core.mem_do_prefetch ),
    .S(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__and2_1 _20860_ (.A(_10317_),
    .B(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _20861_ (.A(_04312_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_2 _20862_ (.A(_06010_),
    .X(_04313_));
 sky130_fd_sc_hd__a21bo_1 _20863_ (.A1(\core.reg_out[2] ),
    .A2(_04313_),
    .B1_N(_06624_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _20864_ (.A0(_04314_),
    .A1(_04699_),
    .S(_06059_),
    .X(_04315_));
 sky130_fd_sc_hd__mux2_1 _20865_ (.A0(_04315_),
    .A1(net55),
    .S(_06055_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _20866_ (.A(_04316_),
    .X(_01528_));
 sky130_fd_sc_hd__a21bo_1 _20867_ (.A1(\core.reg_out[3] ),
    .A2(_04313_),
    .B1_N(_06643_),
    .X(_04317_));
 sky130_fd_sc_hd__mux2_1 _20868_ (.A0(_04317_),
    .A1(_04677_),
    .S(_06059_),
    .X(_04318_));
 sky130_fd_sc_hd__mux2_1 _20869_ (.A0(_04318_),
    .A1(net58),
    .S(_06055_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _20870_ (.A(_04319_),
    .X(_01529_));
 sky130_fd_sc_hd__a21bo_1 _20871_ (.A1(\core.reg_out[4] ),
    .A2(_04313_),
    .B1_N(_06671_),
    .X(_04320_));
 sky130_fd_sc_hd__mux2_1 _20872_ (.A0(_04320_),
    .A1(_04723_),
    .S(_06059_),
    .X(_04321_));
 sky130_fd_sc_hd__mux2_1 _20873_ (.A0(_04321_),
    .A1(net59),
    .S(_06055_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _20874_ (.A(_04322_),
    .X(_01530_));
 sky130_fd_sc_hd__a21bo_1 _20875_ (.A1(\core.reg_out[5] ),
    .A2(_04313_),
    .B1_N(_06697_),
    .X(_04323_));
 sky130_fd_sc_hd__mux2_1 _20876_ (.A0(_04323_),
    .A1(_04728_),
    .S(_06059_),
    .X(_04324_));
 sky130_fd_sc_hd__mux2_1 _20877_ (.A0(_04324_),
    .A1(net60),
    .S(_06055_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _20878_ (.A(_04325_),
    .X(_01531_));
 sky130_fd_sc_hd__a21bo_1 _20879_ (.A1(\core.reg_out[6] ),
    .A2(_04313_),
    .B1_N(_06717_),
    .X(_04326_));
 sky130_fd_sc_hd__mux2_1 _20880_ (.A0(_04326_),
    .A1(_04737_),
    .S(_06059_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_2 _20881_ (.A(_05972_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_1 _20882_ (.A0(_04327_),
    .A1(net61),
    .S(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _20883_ (.A(_04329_),
    .X(_01532_));
 sky130_fd_sc_hd__a21bo_1 _20884_ (.A1(\core.reg_out[7] ),
    .A2(_04313_),
    .B1_N(_06736_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_1 _20885_ (.A0(_04330_),
    .A1(_04734_),
    .S(_05952_),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _20886_ (.A0(_04331_),
    .A1(net62),
    .S(_04328_),
    .X(_04332_));
 sky130_fd_sc_hd__buf_1 _20887_ (.A(_04332_),
    .X(_01533_));
 sky130_fd_sc_hd__clkbuf_2 _20888_ (.A(_05953_),
    .X(_04333_));
 sky130_fd_sc_hd__o211a_1 _20889_ (.A1(_06755_),
    .A2(_05990_),
    .B1(_05982_),
    .C1(_06759_),
    .X(_04334_));
 sky130_fd_sc_hd__a21oi_1 _20890_ (.A1(_04783_),
    .A2(_04333_),
    .B1(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__mux2_1 _20891_ (.A0(_04335_),
    .A1(net63),
    .S(_04328_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _20892_ (.A(_04336_),
    .X(_01534_));
 sky130_fd_sc_hd__a21bo_1 _20893_ (.A1(\core.reg_out[9] ),
    .A2(_06010_),
    .B1_N(_06780_),
    .X(_04337_));
 sky130_fd_sc_hd__mux2_1 _20894_ (.A0(_04337_),
    .A1(_04752_),
    .S(_05952_),
    .X(_04338_));
 sky130_fd_sc_hd__mux2_1 _20895_ (.A0(_04338_),
    .A1(net64),
    .S(_04328_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _20896_ (.A(_04339_),
    .X(_01535_));
 sky130_fd_sc_hd__o211a_1 _20897_ (.A1(_06805_),
    .A2(_05990_),
    .B1(_05982_),
    .C1(_06809_),
    .X(_04340_));
 sky130_fd_sc_hd__a21oi_1 _20898_ (.A1(_04790_),
    .A2(_04333_),
    .B1(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__mux2_1 _20899_ (.A0(_04341_),
    .A1(net35),
    .S(_04328_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _20900_ (.A(_04342_),
    .X(_01536_));
 sky130_fd_sc_hd__clkbuf_2 _20901_ (.A(_05960_),
    .X(_04343_));
 sky130_fd_sc_hd__o211a_1 _20902_ (.A1(_06827_),
    .A2(_05990_),
    .B1(_04343_),
    .C1(_06831_),
    .X(_04344_));
 sky130_fd_sc_hd__a21oi_1 _20903_ (.A1(_04792_),
    .A2(_04333_),
    .B1(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__mux2_1 _20904_ (.A0(_04345_),
    .A1(net36),
    .S(_04328_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _20905_ (.A(_04346_),
    .X(_01537_));
 sky130_fd_sc_hd__o211a_1 _20906_ (.A1(_06852_),
    .A2(_05989_),
    .B1(_04343_),
    .C1(_06856_),
    .X(_04347_));
 sky130_fd_sc_hd__a21oi_1 _20907_ (.A1(_04796_),
    .A2(_04333_),
    .B1(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__mux2_1 _20908_ (.A0(_04348_),
    .A1(net37),
    .S(_09945_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _20909_ (.A(_04349_),
    .X(_01538_));
 sky130_fd_sc_hd__o211a_1 _20910_ (.A1(_06876_),
    .A2(_05989_),
    .B1(_04343_),
    .C1(_06880_),
    .X(_04350_));
 sky130_fd_sc_hd__a21oi_1 _20911_ (.A1(_04799_),
    .A2(_04333_),
    .B1(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__mux2_1 _20912_ (.A0(_04351_),
    .A1(net38),
    .S(_09945_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _20913_ (.A(_04352_),
    .X(_01539_));
 sky130_fd_sc_hd__o211a_1 _20914_ (.A1(_06905_),
    .A2(_05989_),
    .B1(_04343_),
    .C1(_06909_),
    .X(_04353_));
 sky130_fd_sc_hd__a21oi_1 _20915_ (.A1(_04804_),
    .A2(_04333_),
    .B1(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__mux2_1 _20916_ (.A0(_04354_),
    .A1(net39),
    .S(_09945_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _20917_ (.A(_04355_),
    .X(_01540_));
 sky130_fd_sc_hd__o211a_1 _20918_ (.A1(_06928_),
    .A2(_05989_),
    .B1(_04343_),
    .C1(_06932_),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_1 _20919_ (.A1(_04806_),
    .A2(_05953_),
    .B1(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__mux2_1 _20920_ (.A0(_04357_),
    .A1(net40),
    .S(_09945_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _20921_ (.A(_04358_),
    .X(_01541_));
 sky130_fd_sc_hd__o211a_1 _20922_ (.A1(_06960_),
    .A2(_05989_),
    .B1(_04343_),
    .C1(_06964_),
    .X(_04359_));
 sky130_fd_sc_hd__a21oi_1 _20923_ (.A1(_04901_),
    .A2(_05953_),
    .B1(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__mux2_1 _20924_ (.A0(_04360_),
    .A1(net41),
    .S(_09945_),
    .X(_04361_));
 sky130_fd_sc_hd__buf_1 _20925_ (.A(_04361_),
    .X(_01542_));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(clknet_leaf_31_clk),
    .D(_00037_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00038_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _20928_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00039_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _20929_ (.CLK(clknet_3_4__leaf_clk),
    .D(_00040_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_60_clk),
    .D(_00041_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_54_clk),
    .D(_00042_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_27_clk),
    .D(_00043_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_2 _20933_ (.CLK(clknet_leaf_10_clk),
    .D(_00044_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_12_clk),
    .D(_00045_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_2 _20935_ (.CLK(clknet_leaf_29_clk),
    .D(_00046_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_27_clk),
    .D(_00047_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_56_clk),
    .D(_00048_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_7_clk),
    .D(_00049_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(clknet_leaf_92_clk),
    .D(_00050_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(clknet_leaf_58_clk),
    .D(_00051_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _20941_ (.CLK(clknet_leaf_21_clk),
    .D(_01543_),
    .Q(\core.reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20942_ (.CLK(clknet_leaf_21_clk),
    .D(_01554_),
    .Q(\core.reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20943_ (.CLK(clknet_leaf_3_clk),
    .D(_01565_),
    .Q(\core.reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20944_ (.CLK(clknet_leaf_22_clk),
    .D(_01568_),
    .Q(\core.reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_5_clk),
    .D(_01569_),
    .Q(\core.reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20946_ (.CLK(clknet_leaf_3_clk),
    .D(_01570_),
    .Q(\core.reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_4_clk),
    .D(_01571_),
    .Q(\core.reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20948_ (.CLK(clknet_leaf_18_clk),
    .D(_01572_),
    .Q(\core.reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_5_clk),
    .D(_01573_),
    .Q(\core.reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20950_ (.CLK(clknet_leaf_5_clk),
    .D(_01574_),
    .Q(\core.reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20951_ (.CLK(clknet_leaf_20_clk),
    .D(_01544_),
    .Q(\core.reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20952_ (.CLK(clknet_leaf_6_clk),
    .D(_01545_),
    .Q(\core.reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20953_ (.CLK(clknet_leaf_19_clk),
    .D(_01546_),
    .Q(\core.reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20954_ (.CLK(clknet_leaf_19_clk),
    .D(_01547_),
    .Q(\core.reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(clknet_leaf_20_clk),
    .D(_01548_),
    .Q(\core.reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20956_ (.CLK(clknet_leaf_5_clk),
    .D(_01549_),
    .Q(\core.reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(clknet_leaf_6_clk),
    .D(_01550_),
    .Q(\core.reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20958_ (.CLK(clknet_leaf_26_clk),
    .D(_01551_),
    .Q(\core.reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20959_ (.CLK(clknet_leaf_20_clk),
    .D(_01552_),
    .Q(\core.reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20960_ (.CLK(clknet_leaf_20_clk),
    .D(_01553_),
    .Q(\core.reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20961_ (.CLK(clknet_leaf_25_clk),
    .D(_01555_),
    .Q(\core.reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(clknet_leaf_18_clk),
    .D(_01556_),
    .Q(\core.reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20963_ (.CLK(clknet_leaf_20_clk),
    .D(_01557_),
    .Q(\core.reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(clknet_leaf_20_clk),
    .D(_01558_),
    .Q(\core.reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_19_clk),
    .D(_01559_),
    .Q(\core.reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20966_ (.CLK(clknet_leaf_19_clk),
    .D(_01560_),
    .Q(\core.reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(clknet_leaf_25_clk),
    .D(_01561_),
    .Q(\core.reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_21_clk),
    .D(_01562_),
    .Q(\core.reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_25_clk),
    .D(_01563_),
    .Q(\core.reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_18_clk),
    .D(_01564_),
    .Q(\core.reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_21_clk),
    .D(_01566_),
    .Q(\core.reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_21_clk),
    .D(_01567_),
    .Q(\core.reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20973_ (.CLK(clknet_leaf_23_clk),
    .D(_00052_),
    .Q(\core.pcpi_rs1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_16_clk),
    .D(_00053_),
    .Q(\core.count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_18_clk),
    .D(_00054_),
    .Q(\core.count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_19_clk),
    .D(_00055_),
    .Q(\core.count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_17_clk),
    .D(_00056_),
    .Q(\core.count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20978_ (.CLK(clknet_leaf_17_clk),
    .D(_00057_),
    .Q(\core.count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_17_clk),
    .D(_00058_),
    .Q(\core.count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_17_clk),
    .D(_00059_),
    .Q(\core.count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_17_clk),
    .D(_00060_),
    .Q(\core.count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_17_clk),
    .D(_00061_),
    .Q(\core.count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_19_clk),
    .D(_00062_),
    .Q(\core.count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20984_ (.CLK(clknet_leaf_16_clk),
    .D(_00063_),
    .Q(\core.count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20985_ (.CLK(clknet_leaf_16_clk),
    .D(_00064_),
    .Q(\core.count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20986_ (.CLK(clknet_leaf_16_clk),
    .D(_00065_),
    .Q(\core.count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20987_ (.CLK(clknet_leaf_16_clk),
    .D(_00066_),
    .Q(\core.count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_17_clk),
    .D(_00067_),
    .Q(\core.count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_13_clk),
    .D(_00068_),
    .Q(\core.count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_16_clk),
    .D(_00069_),
    .Q(\core.count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_20_clk),
    .D(_00070_),
    .Q(\core.count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20992_ (.CLK(clknet_leaf_13_clk),
    .D(_00071_),
    .Q(\core.count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_17_clk),
    .D(_00072_),
    .Q(\core.count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_16_clk),
    .D(_00073_),
    .Q(\core.count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_15_clk),
    .D(_00074_),
    .Q(\core.count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_13_clk),
    .D(_00075_),
    .Q(\core.count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_leaf_13_clk),
    .D(_00076_),
    .Q(\core.count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20998_ (.CLK(clknet_leaf_13_clk),
    .D(_00077_),
    .Q(\core.count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20999_ (.CLK(clknet_leaf_14_clk),
    .D(_00078_),
    .Q(\core.count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_20_clk),
    .D(_00079_),
    .Q(\core.count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_2 _21001_ (.CLK(clknet_leaf_15_clk),
    .D(_00080_),
    .Q(\core.count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_15_clk),
    .D(_00081_),
    .Q(\core.count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _21003_ (.CLK(clknet_leaf_13_clk),
    .D(_00082_),
    .Q(\core.count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_15_clk),
    .D(_00083_),
    .Q(\core.count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _21005_ (.CLK(clknet_leaf_14_clk),
    .D(_00084_),
    .Q(\core.count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_14_clk),
    .D(_00085_),
    .Q(\core.count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21007_ (.CLK(clknet_leaf_15_clk),
    .D(_00086_),
    .Q(\core.count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_16_clk),
    .D(_00087_),
    .Q(\core.count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21009_ (.CLK(clknet_leaf_16_clk),
    .D(_00088_),
    .Q(\core.count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_2 _21010_ (.CLK(clknet_leaf_15_clk),
    .D(_00089_),
    .Q(\core.count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_2 _21011_ (.CLK(clknet_leaf_15_clk),
    .D(_00090_),
    .Q(\core.count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21012_ (.CLK(clknet_leaf_15_clk),
    .D(_00091_),
    .Q(\core.count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21013_ (.CLK(clknet_leaf_16_clk),
    .D(_00092_),
    .Q(\core.count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_2 _21014_ (.CLK(clknet_leaf_16_clk),
    .D(_00093_),
    .Q(\core.count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_15_clk),
    .D(_00094_),
    .Q(\core.count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_2 _21016_ (.CLK(clknet_leaf_16_clk),
    .D(_00095_),
    .Q(\core.count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_16_clk),
    .D(_00096_),
    .Q(\core.count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_14_clk),
    .D(_00097_),
    .Q(\core.count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00098_),
    .Q(\core.count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_2 _21020_ (.CLK(clknet_leaf_14_clk),
    .D(_00099_),
    .Q(\core.count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_15_clk),
    .D(_00100_),
    .Q(\core.count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_2 _21022_ (.CLK(clknet_leaf_15_clk),
    .D(_00101_),
    .Q(\core.count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_15_clk),
    .D(_00102_),
    .Q(\core.count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_14_clk),
    .D(_00103_),
    .Q(\core.count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(clknet_leaf_16_clk),
    .D(_00104_),
    .Q(\core.count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_14_clk),
    .D(_00105_),
    .Q(\core.count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 _21027_ (.CLK(clknet_leaf_14_clk),
    .D(_00106_),
    .Q(\core.count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_14_clk),
    .D(_00107_),
    .Q(\core.count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21029_ (.CLK(clknet_leaf_15_clk),
    .D(_00108_),
    .Q(\core.count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_14_clk),
    .D(_00109_),
    .Q(\core.count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_2 _21031_ (.CLK(clknet_leaf_13_clk),
    .D(_00110_),
    .Q(\core.count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_2 _21032_ (.CLK(clknet_leaf_13_clk),
    .D(_00111_),
    .Q(\core.count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_15_clk),
    .D(_00112_),
    .Q(\core.count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_2 _21034_ (.CLK(clknet_leaf_14_clk),
    .D(_00113_),
    .Q(\core.count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_14_clk),
    .D(_00114_),
    .Q(\core.count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_15_clk),
    .D(_00115_),
    .Q(\core.count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(clknet_leaf_15_clk),
    .D(_00116_),
    .Q(\core.count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_18_clk),
    .D(_00117_),
    .Q(\core.reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(clknet_leaf_5_clk),
    .D(_00118_),
    .Q(\core.reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_5_clk),
    .D(_00119_),
    .Q(\core.reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_4 _21041_ (.CLK(clknet_leaf_6_clk),
    .D(_00120_),
    .Q(\core.reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_5_clk),
    .D(_00121_),
    .Q(\core.reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(clknet_leaf_17_clk),
    .D(_00122_),
    .Q(\core.reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_5_clk),
    .D(_00123_),
    .Q(\core.reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_6_clk),
    .D(_00124_),
    .Q(\core.reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21046_ (.CLK(clknet_leaf_6_clk),
    .D(_00125_),
    .Q(\core.reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21047_ (.CLK(clknet_leaf_19_clk),
    .D(_00126_),
    .Q(\core.reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_18_clk),
    .D(_00127_),
    .Q(\core.reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_17_clk),
    .D(_00128_),
    .Q(\core.reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(clknet_leaf_18_clk),
    .D(net136),
    .Q(\core.reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_25_clk),
    .D(_00130_),
    .Q(\core.reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(clknet_leaf_18_clk),
    .D(_00131_),
    .Q(\core.reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21053_ (.CLK(clknet_leaf_17_clk),
    .D(_00132_),
    .Q(\core.reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21054_ (.CLK(clknet_leaf_20_clk),
    .D(_00133_),
    .Q(\core.reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_5_clk),
    .D(_00134_),
    .Q(\core.reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_5_clk),
    .D(_00135_),
    .Q(\core.reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_26_clk),
    .D(_00136_),
    .Q(\core.reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_leaf_25_clk),
    .D(_00137_),
    .Q(\core.reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_20_clk),
    .D(_00138_),
    .Q(\core.reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(clknet_leaf_20_clk),
    .D(_00139_),
    .Q(\core.reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(clknet_leaf_26_clk),
    .D(_00140_),
    .Q(\core.reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(clknet_leaf_26_clk),
    .D(_00141_),
    .Q(\core.reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_20_clk),
    .D(_00142_),
    .Q(\core.reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_20_clk),
    .D(_00143_),
    .Q(\core.reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_26_clk),
    .D(_00144_),
    .Q(\core.reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_19_clk),
    .D(_00145_),
    .Q(\core.reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_18_clk),
    .D(_00146_),
    .Q(\core.reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(clknet_leaf_18_clk),
    .D(_00147_),
    .Q(\core.reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_3_clk),
    .D(_00148_),
    .Q(\core.reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_3_clk),
    .D(_00149_),
    .Q(\core.reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21071_ (.CLK(clknet_leaf_3_clk),
    .D(_00150_),
    .Q(\core.reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_0_clk),
    .D(_00151_),
    .Q(\core.reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21073_ (.CLK(clknet_leaf_3_clk),
    .D(_00152_),
    .Q(\core.reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21074_ (.CLK(clknet_leaf_1_clk),
    .D(_00153_),
    .Q(\core.reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_0_clk),
    .D(_00154_),
    .Q(\core.reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_21_clk),
    .D(_00155_),
    .Q(\core.reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_21_clk),
    .D(_00156_),
    .Q(\core.reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_22_clk),
    .D(_00157_),
    .Q(\core.reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_3_clk),
    .D(_00158_),
    .Q(\core.reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(clknet_leaf_3_clk),
    .D(_00159_),
    .Q(\core.reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(clknet_leaf_22_clk),
    .D(_00160_),
    .Q(\core.reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_2_clk),
    .D(_00161_),
    .Q(\core.reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_23_clk),
    .D(_00162_),
    .Q(\core.reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_22_clk),
    .D(_00163_),
    .Q(\core.reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_23_clk),
    .D(_00164_),
    .Q(\core.reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_24_clk),
    .D(_00165_),
    .Q(\core.reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_21_clk),
    .D(_00166_),
    .Q(\core.reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _21088_ (.CLK(clknet_leaf_25_clk),
    .D(_00167_),
    .Q(\core.reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_24_clk),
    .D(_00168_),
    .Q(\core.reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_24_clk),
    .D(_00169_),
    .Q(\core.reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(clknet_leaf_24_clk),
    .D(_00170_),
    .Q(\core.reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_4 _21092_ (.CLK(clknet_leaf_25_clk),
    .D(_00171_),
    .Q(\core.reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_4 _21093_ (.CLK(clknet_leaf_25_clk),
    .D(_00172_),
    .Q(\core.reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_21_clk),
    .D(_00173_),
    .Q(\core.reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_23_clk),
    .D(_00174_),
    .Q(\core.reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_23_clk),
    .D(_00175_),
    .Q(\core.reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _21097_ (.CLK(clknet_leaf_24_clk),
    .D(_00176_),
    .Q(\core.reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(clknet_leaf_23_clk),
    .D(_00177_),
    .Q(\core.reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _21099_ (.CLK(clknet_leaf_24_clk),
    .D(_00178_),
    .Q(\core.reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(clknet_leaf_16_clk),
    .D(_00179_),
    .Q(\core.count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(clknet_leaf_14_clk),
    .D(_00180_),
    .Q(\core.count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(clknet_leaf_16_clk),
    .D(_00181_),
    .Q(\core.count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(clknet_leaf_14_clk),
    .D(_00182_),
    .Q(\core.count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21104_ (.CLK(clknet_leaf_15_clk),
    .D(_00183_),
    .Q(\core.count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(clknet_leaf_16_clk),
    .D(_00184_),
    .Q(\core.count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(clknet_leaf_15_clk),
    .D(_00185_),
    .Q(\core.count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(clknet_leaf_15_clk),
    .D(_00186_),
    .Q(\core.count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(clknet_leaf_16_clk),
    .D(_00187_),
    .Q(\core.count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(clknet_leaf_16_clk),
    .D(_00188_),
    .Q(\core.count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(clknet_leaf_16_clk),
    .D(_00189_),
    .Q(\core.count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(clknet_leaf_14_clk),
    .D(_00190_),
    .Q(\core.count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(clknet_leaf_15_clk),
    .D(_00191_),
    .Q(\core.count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21113_ (.CLK(clknet_leaf_15_clk),
    .D(_00192_),
    .Q(\core.count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(clknet_leaf_14_clk),
    .D(_00193_),
    .Q(\core.count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(clknet_leaf_14_clk),
    .D(_00194_),
    .Q(\core.count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(clknet_leaf_14_clk),
    .D(_00195_),
    .Q(\core.count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(clknet_leaf_14_clk),
    .D(_00196_),
    .Q(\core.count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(clknet_leaf_13_clk),
    .D(_00197_),
    .Q(\core.count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(clknet_leaf_13_clk),
    .D(_00198_),
    .Q(\core.count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(clknet_leaf_13_clk),
    .D(_00199_),
    .Q(\core.count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_14_clk),
    .D(_00200_),
    .Q(\core.count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(clknet_leaf_13_clk),
    .D(_00201_),
    .Q(\core.count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_13_clk),
    .D(_00202_),
    .Q(\core.count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_14_clk),
    .D(_00203_),
    .Q(\core.count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _21125_ (.CLK(clknet_leaf_13_clk),
    .D(_00204_),
    .Q(\core.count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_13_clk),
    .D(_00205_),
    .Q(\core.count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_14_clk),
    .D(_00206_),
    .Q(\core.count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_15_clk),
    .D(_00207_),
    .Q(\core.count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(clknet_leaf_15_clk),
    .D(_00208_),
    .Q(\core.count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _21130_ (.CLK(clknet_leaf_16_clk),
    .D(_00209_),
    .Q(\core.count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_15_clk),
    .D(_00210_),
    .Q(\core.count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_20_clk),
    .D(_00211_),
    .Q(\core.count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_2 _21133_ (.CLK(clknet_leaf_13_clk),
    .D(_00212_),
    .Q(\core.count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_16_clk),
    .D(_00213_),
    .Q(\core.count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_16_clk),
    .D(_00214_),
    .Q(\core.count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_2 _21136_ (.CLK(clknet_leaf_16_clk),
    .D(_00215_),
    .Q(\core.count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_15_clk),
    .D(_00216_),
    .Q(\core.count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21138_ (.CLK(clknet_leaf_16_clk),
    .D(_00217_),
    .Q(\core.count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21139_ (.CLK(clknet_leaf_14_clk),
    .D(_00218_),
    .Q(\core.count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_2 _21140_ (.CLK(clknet_leaf_17_clk),
    .D(_00219_),
    .Q(\core.count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_2 _21141_ (.CLK(clknet_leaf_19_clk),
    .D(_00220_),
    .Q(\core.count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21142_ (.CLK(clknet_leaf_13_clk),
    .D(_00221_),
    .Q(\core.count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21143_ (.CLK(clknet_leaf_20_clk),
    .D(_00222_),
    .Q(\core.count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21144_ (.CLK(clknet_leaf_19_clk),
    .D(_00223_),
    .Q(\core.count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21145_ (.CLK(clknet_leaf_13_clk),
    .D(_00224_),
    .Q(\core.count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21146_ (.CLK(clknet_leaf_14_clk),
    .D(_00225_),
    .Q(\core.count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21147_ (.CLK(clknet_leaf_19_clk),
    .D(_00226_),
    .Q(\core.count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21148_ (.CLK(clknet_leaf_19_clk),
    .D(_00227_),
    .Q(\core.count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_2 _21149_ (.CLK(clknet_leaf_19_clk),
    .D(_00228_),
    .Q(\core.count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(clknet_leaf_19_clk),
    .D(_00229_),
    .Q(\core.count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21151_ (.CLK(clknet_leaf_19_clk),
    .D(_00230_),
    .Q(\core.count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(clknet_leaf_19_clk),
    .D(_00231_),
    .Q(\core.count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21153_ (.CLK(clknet_leaf_13_clk),
    .D(_00232_),
    .Q(\core.count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_13_clk),
    .D(_00233_),
    .Q(\core.count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(clknet_leaf_13_clk),
    .D(_00234_),
    .Q(\core.count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_2 _21156_ (.CLK(clknet_leaf_13_clk),
    .D(_00235_),
    .Q(\core.count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_14_clk),
    .D(_00236_),
    .Q(\core.count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(clknet_leaf_13_clk),
    .D(_00237_),
    .Q(\core.count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_2 _21159_ (.CLK(clknet_leaf_20_clk),
    .D(_00238_),
    .Q(\core.count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_13_clk),
    .D(_00239_),
    .Q(\core.count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_20_clk),
    .D(_00240_),
    .Q(\core.count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_2 _21162_ (.CLK(clknet_leaf_13_clk),
    .D(_00241_),
    .Q(\core.count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_2 _21163_ (.CLK(clknet_leaf_19_clk),
    .D(_00242_),
    .Q(\core.count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_2_clk),
    .D(_00243_),
    .Q(\core.pcpi_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_1_clk),
    .D(_00244_),
    .Q(\core.pcpi_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(clknet_leaf_1_clk),
    .D(_00245_),
    .Q(\core.pcpi_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_0_clk),
    .D(_00246_),
    .Q(\core.pcpi_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_4_clk),
    .D(_00247_),
    .Q(\core.pcpi_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_0_clk),
    .D(_00248_),
    .Q(\core.pcpi_rs1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_2_clk),
    .D(_00249_),
    .Q(\core.pcpi_rs1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_0_clk),
    .D(_00250_),
    .Q(\core.pcpi_rs1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_0_clk),
    .D(_00251_),
    .Q(\core.pcpi_rs1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_0_clk),
    .D(_00252_),
    .Q(\core.pcpi_rs1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_2_clk),
    .D(_00253_),
    .Q(\core.pcpi_rs1[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21175_ (.CLK(clknet_leaf_1_clk),
    .D(_00254_),
    .Q(\core.pcpi_rs1[11] ));
 sky130_fd_sc_hd__dfxtp_4 _21176_ (.CLK(clknet_leaf_23_clk),
    .D(_00255_),
    .Q(\core.pcpi_rs1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21177_ (.CLK(clknet_leaf_1_clk),
    .D(_00256_),
    .Q(\core.pcpi_rs1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_23_clk),
    .D(_00257_),
    .Q(\core.pcpi_rs1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_1_clk),
    .D(_00258_),
    .Q(\core.pcpi_rs1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_1_clk),
    .D(_00259_),
    .Q(\core.pcpi_rs1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_23_clk),
    .D(_00260_),
    .Q(\core.pcpi_rs1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _21182_ (.CLK(clknet_leaf_23_clk),
    .D(_00261_),
    .Q(\core.pcpi_rs1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_1_clk),
    .D(_00262_),
    .Q(\core.pcpi_rs1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _21184_ (.CLK(clknet_leaf_23_clk),
    .D(_00263_),
    .Q(\core.pcpi_rs1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_1_clk),
    .D(_00264_),
    .Q(\core.pcpi_rs1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_1_clk),
    .D(_00265_),
    .Q(\core.pcpi_rs1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_2_clk),
    .D(_00266_),
    .Q(\core.pcpi_rs1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_1_clk),
    .D(_00267_),
    .Q(\core.pcpi_rs1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _21189_ (.CLK(clknet_leaf_23_clk),
    .D(_00268_),
    .Q(\core.pcpi_rs1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_23_clk),
    .D(_00269_),
    .Q(\core.pcpi_rs1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_1_clk),
    .D(_00270_),
    .Q(\core.pcpi_rs1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_23_clk),
    .D(_00271_),
    .Q(\core.pcpi_rs1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_1_clk),
    .D(_00272_),
    .Q(\core.pcpi_rs1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_1_clk),
    .D(_00273_),
    .Q(\core.pcpi_rs1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _21195_ (.CLK(clknet_leaf_36_clk),
    .D(_00274_),
    .Q(\core.mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21196_ (.CLK(clknet_leaf_36_clk),
    .D(_00275_),
    .Q(\core.mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_70_clk),
    .D(_00276_),
    .Q(\core.cpuregs[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 _21198_ (.CLK(clknet_leaf_68_clk),
    .D(_00277_),
    .Q(\core.cpuregs[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_84_clk),
    .D(_00278_),
    .Q(\core.cpuregs[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_84_clk),
    .D(_00279_),
    .Q(\core.cpuregs[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_67_clk),
    .D(_00280_),
    .Q(\core.cpuregs[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_74_clk),
    .D(_00281_),
    .Q(\core.cpuregs[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_74_clk),
    .D(_00282_),
    .Q(\core.cpuregs[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_67_clk),
    .D(_00283_),
    .Q(\core.cpuregs[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_67_clk),
    .D(_00284_),
    .Q(\core.cpuregs[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 _21206_ (.CLK(clknet_leaf_67_clk),
    .D(_00285_),
    .Q(\core.cpuregs[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_68_clk),
    .D(_00286_),
    .Q(\core.cpuregs[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_56_clk),
    .D(_00287_),
    .Q(\core.cpuregs[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_44_clk),
    .D(_00288_),
    .Q(\core.cpuregs[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 _21210_ (.CLK(clknet_leaf_44_clk),
    .D(_00289_),
    .Q(\core.cpuregs[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_44_clk),
    .D(_00290_),
    .Q(\core.cpuregs[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(clknet_leaf_71_clk),
    .D(_00291_),
    .Q(\core.cpuregs[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_72_clk),
    .D(_00292_),
    .Q(\core.cpuregs[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_44_clk),
    .D(_00293_),
    .Q(\core.cpuregs[23][17] ));
 sky130_fd_sc_hd__dfxtp_2 _21215_ (.CLK(clknet_leaf_71_clk),
    .D(_00294_),
    .Q(\core.cpuregs[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_62_clk),
    .D(_00295_),
    .Q(\core.cpuregs[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_61_clk),
    .D(_00296_),
    .Q(\core.cpuregs[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_55_clk),
    .D(_00297_),
    .Q(\core.cpuregs[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_62_clk),
    .D(_00298_),
    .Q(\core.cpuregs[23][22] ));
 sky130_fd_sc_hd__dfxtp_2 _21220_ (.CLK(clknet_leaf_54_clk),
    .D(_00299_),
    .Q(\core.cpuregs[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_54_clk),
    .D(_00300_),
    .Q(\core.cpuregs[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_62_clk),
    .D(_00301_),
    .Q(\core.cpuregs[23][25] ));
 sky130_fd_sc_hd__dfxtp_4 _21223_ (.CLK(clknet_leaf_69_clk),
    .D(_00302_),
    .Q(\core.cpuregs[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_55_clk),
    .D(_00303_),
    .Q(\core.cpuregs[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_69_clk),
    .D(_00304_),
    .Q(\core.cpuregs[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_62_clk),
    .D(_00305_),
    .Q(\core.cpuregs[23][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21227_ (.CLK(clknet_leaf_63_clk),
    .D(_00306_),
    .Q(\core.cpuregs[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_70_clk),
    .D(_00307_),
    .Q(\core.cpuregs[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_70_clk),
    .D(_00308_),
    .Q(\core.cpuregs[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_70_clk),
    .D(_00309_),
    .Q(\core.cpuregs[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_67_clk),
    .D(_00310_),
    .Q(\core.cpuregs[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_84_clk),
    .D(_00311_),
    .Q(\core.cpuregs[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_83_clk),
    .D(_00312_),
    .Q(\core.cpuregs[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_67_clk),
    .D(_00313_),
    .Q(\core.cpuregs[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_67_clk),
    .D(_00314_),
    .Q(\core.cpuregs[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_67_clk),
    .D(_00315_),
    .Q(\core.cpuregs[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_68_clk),
    .D(_00316_),
    .Q(\core.cpuregs[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_71_clk),
    .D(_00317_),
    .Q(\core.cpuregs[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_68_clk),
    .D(_00318_),
    .Q(\core.cpuregs[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_45_clk),
    .D(_00319_),
    .Q(\core.cpuregs[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_72_clk),
    .D(_00320_),
    .Q(\core.cpuregs[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_56_clk),
    .D(_00321_),
    .Q(\core.cpuregs[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_43_clk),
    .D(_00322_),
    .Q(\core.cpuregs[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_43_clk),
    .D(_00323_),
    .Q(\core.cpuregs[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_72_clk),
    .D(_00324_),
    .Q(\core.cpuregs[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_44_clk),
    .D(_00325_),
    .Q(\core.cpuregs[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(clknet_leaf_56_clk),
    .D(_00326_),
    .Q(\core.cpuregs[30][18] ));
 sky130_fd_sc_hd__dfxtp_2 _21248_ (.CLK(clknet_leaf_52_clk),
    .D(_00327_),
    .Q(\core.cpuregs[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_53_clk),
    .D(_00328_),
    .Q(\core.cpuregs[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_56_clk),
    .D(_00329_),
    .Q(\core.cpuregs[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_55_clk),
    .D(_00330_),
    .Q(\core.cpuregs[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_53_clk),
    .D(_00331_),
    .Q(\core.cpuregs[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_55_clk),
    .D(_00332_),
    .Q(\core.cpuregs[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_56_clk),
    .D(_00333_),
    .Q(\core.cpuregs[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_62_clk),
    .D(_00334_),
    .Q(\core.cpuregs[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_58_clk),
    .D(_00335_),
    .Q(\core.cpuregs[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_57_clk),
    .D(_00336_),
    .Q(\core.cpuregs[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_69_clk),
    .D(_00337_),
    .Q(\core.cpuregs[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_58_clk),
    .D(_00338_),
    .Q(\core.cpuregs[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_69_clk),
    .D(_00339_),
    .Q(\core.cpuregs[30][31] ));
 sky130_fd_sc_hd__dfxtp_2 _21261_ (.CLK(clknet_leaf_2_clk),
    .D(_00340_),
    .Q(\core.reg_sh[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_22_clk),
    .D(_00341_),
    .Q(\core.reg_sh[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_71_clk),
    .D(_00342_),
    .Q(\core.cpuregs[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_45_clk),
    .D(_00343_),
    .Q(\core.cpuregs[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_85_clk),
    .D(_00344_),
    .Q(\core.cpuregs[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_84_clk),
    .D(_00345_),
    .Q(\core.cpuregs[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_85_clk),
    .D(_00346_),
    .Q(\core.cpuregs[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_67_clk),
    .D(_00347_),
    .Q(\core.cpuregs[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_72_clk),
    .D(_00348_),
    .Q(\core.cpuregs[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_82_clk),
    .D(_00349_),
    .Q(\core.cpuregs[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_67_clk),
    .D(_00350_),
    .Q(\core.cpuregs[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_68_clk),
    .D(_00351_),
    .Q(\core.cpuregs[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_67_clk),
    .D(_00352_),
    .Q(\core.cpuregs[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_56_clk),
    .D(_00353_),
    .Q(\core.cpuregs[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_69_clk),
    .D(_00354_),
    .Q(\core.cpuregs[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 _21276_ (.CLK(clknet_leaf_71_clk),
    .D(_00355_),
    .Q(\core.cpuregs[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21277_ (.CLK(clknet_leaf_44_clk),
    .D(_00356_),
    .Q(\core.cpuregs[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21278_ (.CLK(clknet_leaf_72_clk),
    .D(_00357_),
    .Q(\core.cpuregs[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_72_clk),
    .D(_00358_),
    .Q(\core.cpuregs[22][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21280_ (.CLK(clknet_leaf_45_clk),
    .D(_00359_),
    .Q(\core.cpuregs[22][17] ));
 sky130_fd_sc_hd__dfxtp_2 _21281_ (.CLK(clknet_leaf_71_clk),
    .D(_00360_),
    .Q(\core.cpuregs[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_53_clk),
    .D(_00361_),
    .Q(\core.cpuregs[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_53_clk),
    .D(_00362_),
    .Q(\core.cpuregs[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_61_clk),
    .D(_00363_),
    .Q(\core.cpuregs[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_55_clk),
    .D(_00364_),
    .Q(\core.cpuregs[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_53_clk),
    .D(_00365_),
    .Q(\core.cpuregs[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_57_clk),
    .D(_00366_),
    .Q(\core.cpuregs[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_54_clk),
    .D(_00367_),
    .Q(\core.cpuregs[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_57_clk),
    .D(_00368_),
    .Q(\core.cpuregs[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_61_clk),
    .D(_00369_),
    .Q(\core.cpuregs[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_56_clk),
    .D(_00370_),
    .Q(\core.cpuregs[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_57_clk),
    .D(_00371_),
    .Q(\core.cpuregs[22][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21293_ (.CLK(clknet_leaf_69_clk),
    .D(_00372_),
    .Q(\core.cpuregs[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(clknet_leaf_69_clk),
    .D(_00373_),
    .Q(\core.cpuregs[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_44_clk),
    .D(_00374_),
    .Q(\core.cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_46_clk),
    .D(_00375_),
    .Q(\core.cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(clknet_leaf_85_clk),
    .D(_00376_),
    .Q(\core.cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_82_clk),
    .D(_00377_),
    .Q(\core.cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_82_clk),
    .D(_00378_),
    .Q(\core.cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_75_clk),
    .D(_00379_),
    .Q(\core.cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _21301_ (.CLK(clknet_leaf_75_clk),
    .D(_00380_),
    .Q(\core.cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_74_clk),
    .D(_00381_),
    .Q(\core.cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_72_clk),
    .D(_00382_),
    .Q(\core.cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_72_clk),
    .D(_00383_),
    .Q(\core.cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_68_clk),
    .D(_00384_),
    .Q(\core.cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_45_clk),
    .D(_00385_),
    .Q(\core.cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_72_clk),
    .D(_00386_),
    .Q(\core.cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_79_clk),
    .D(_00387_),
    .Q(\core.cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21309_ (.CLK(clknet_leaf_42_clk),
    .D(_00388_),
    .Q(\core.cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21310_ (.CLK(clknet_leaf_45_clk),
    .D(_00389_),
    .Q(\core.cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_43_clk),
    .D(_00390_),
    .Q(\core.cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21312_ (.CLK(clknet_leaf_43_clk),
    .D(_00391_),
    .Q(\core.cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_46_clk),
    .D(_00392_),
    .Q(\core.cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_52_clk),
    .D(_00393_),
    .Q(\core.cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_61_clk),
    .D(_00394_),
    .Q(\core.cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_35_clk),
    .D(_00395_),
    .Q(\core.cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_52_clk),
    .D(_00396_),
    .Q(\core.cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_51_clk),
    .D(_00397_),
    .Q(\core.cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_52_clk),
    .D(_00398_),
    .Q(\core.cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_57_clk),
    .D(_00399_),
    .Q(\core.cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_56_clk),
    .D(_00400_),
    .Q(\core.cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_61_clk),
    .D(_00401_),
    .Q(\core.cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_69_clk),
    .D(_00402_),
    .Q(\core.cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_56_clk),
    .D(_00403_),
    .Q(\core.cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_62_clk),
    .D(_00404_),
    .Q(\core.cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_56_clk),
    .D(_00405_),
    .Q(\core.cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_71_clk),
    .D(_00406_),
    .Q(\core.cpuregs[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _21328_ (.CLK(clknet_leaf_45_clk),
    .D(_00407_),
    .Q(\core.cpuregs[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_67_clk),
    .D(_00408_),
    .Q(\core.cpuregs[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_85_clk),
    .D(_00409_),
    .Q(\core.cpuregs[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_83_clk),
    .D(_00410_),
    .Q(\core.cpuregs[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_67_clk),
    .D(_00411_),
    .Q(\core.cpuregs[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_82_clk),
    .D(_00412_),
    .Q(\core.cpuregs[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_67_clk),
    .D(_00413_),
    .Q(\core.cpuregs[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_71_clk),
    .D(_00414_),
    .Q(\core.cpuregs[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_68_clk),
    .D(_00415_),
    .Q(\core.cpuregs[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_44_clk),
    .D(_00416_),
    .Q(\core.cpuregs[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_45_clk),
    .D(_00417_),
    .Q(\core.cpuregs[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_74_clk),
    .D(_00418_),
    .Q(\core.cpuregs[27][12] ));
 sky130_fd_sc_hd__dfxtp_2 _21340_ (.CLK(clknet_leaf_46_clk),
    .D(_00419_),
    .Q(\core.cpuregs[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_73_clk),
    .D(_00420_),
    .Q(\core.cpuregs[27][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21342_ (.CLK(clknet_leaf_43_clk),
    .D(_00421_),
    .Q(\core.cpuregs[27][15] ));
 sky130_fd_sc_hd__dfxtp_2 _21343_ (.CLK(clknet_leaf_73_clk),
    .D(_00422_),
    .Q(\core.cpuregs[27][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21344_ (.CLK(clknet_leaf_74_clk),
    .D(_00423_),
    .Q(\core.cpuregs[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_71_clk),
    .D(_00424_),
    .Q(\core.cpuregs[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_61_clk),
    .D(_00425_),
    .Q(\core.cpuregs[27][19] ));
 sky130_fd_sc_hd__dfxtp_2 _21347_ (.CLK(clknet_leaf_53_clk),
    .D(_00426_),
    .Q(\core.cpuregs[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_57_clk),
    .D(_00427_),
    .Q(\core.cpuregs[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_53_clk),
    .D(_00428_),
    .Q(\core.cpuregs[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_57_clk),
    .D(_00429_),
    .Q(\core.cpuregs[27][23] ));
 sky130_fd_sc_hd__dfxtp_2 _21351_ (.CLK(clknet_leaf_53_clk),
    .D(_00430_),
    .Q(\core.cpuregs[27][24] ));
 sky130_fd_sc_hd__dfxtp_2 _21352_ (.CLK(clknet_leaf_61_clk),
    .D(_00431_),
    .Q(\core.cpuregs[27][25] ));
 sky130_fd_sc_hd__dfxtp_2 _21353_ (.CLK(clknet_leaf_63_clk),
    .D(_00432_),
    .Q(\core.cpuregs[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_62_clk),
    .D(_00433_),
    .Q(\core.cpuregs[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_61_clk),
    .D(_00434_),
    .Q(\core.cpuregs[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_69_clk),
    .D(_00435_),
    .Q(\core.cpuregs[27][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21357_ (.CLK(clknet_leaf_58_clk),
    .D(_00436_),
    .Q(\core.cpuregs[27][30] ));
 sky130_fd_sc_hd__dfxtp_2 _21358_ (.CLK(clknet_leaf_45_clk),
    .D(_00437_),
    .Q(\core.cpuregs[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_8_clk),
    .D(_00438_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_3_4__leaf_clk),
    .D(_00439_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_60_clk),
    .D(_00440_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_88_clk),
    .D(_00441_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_87_clk),
    .D(_00442_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_86_clk),
    .D(_00443_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_33_clk),
    .D(_00444_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _21366_ (.CLK(clknet_leaf_86_clk),
    .D(_00445_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_91_clk),
    .D(_00446_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_28_clk),
    .D(_00447_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_7_clk),
    .D(_00448_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_91_clk),
    .D(_00449_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_52_clk),
    .D(_00450_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_31_clk),
    .D(_00451_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00452_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_31_clk),
    .D(_00453_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_86_clk),
    .D(_00454_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_10_clk),
    .D(_00455_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_92_clk),
    .D(_00456_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _21378_ (.CLK(clknet_leaf_90_clk),
    .D(_00457_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_10_clk),
    .D(_00458_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_12_clk),
    .D(_00459_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_90_clk),
    .D(_00460_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _21382_ (.CLK(clknet_leaf_10_clk),
    .D(_00461_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _21383_ (.CLK(clknet_leaf_88_clk),
    .D(_00462_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_89_clk),
    .D(_00463_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _21385_ (.CLK(clknet_leaf_29_clk),
    .D(_00464_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_2 _21386_ (.CLK(clknet_leaf_27_clk),
    .D(_00465_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_2 _21387_ (.CLK(clknet_leaf_86_clk),
    .D(_00466_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _21388_ (.CLK(clknet_leaf_29_clk),
    .D(_00467_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_2 _21389_ (.CLK(clknet_leaf_10_clk),
    .D(_00468_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_33_clk),
    .D(_00469_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _21391_ (.CLK(clknet_leaf_29_clk),
    .D(_00470_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_70_clk),
    .D(_00471_),
    .Q(\core.cpuregs[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_44_clk),
    .D(_00472_),
    .Q(\core.cpuregs[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_84_clk),
    .D(_00473_),
    .Q(\core.cpuregs[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_85_clk),
    .D(_00474_),
    .Q(\core.cpuregs[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_85_clk),
    .D(_00475_),
    .Q(\core.cpuregs[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 _21397_ (.CLK(clknet_leaf_74_clk),
    .D(_00476_),
    .Q(\core.cpuregs[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_75_clk),
    .D(_00477_),
    .Q(\core.cpuregs[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_85_clk),
    .D(_00478_),
    .Q(\core.cpuregs[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_68_clk),
    .D(_00479_),
    .Q(\core.cpuregs[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_72_clk),
    .D(_00480_),
    .Q(\core.cpuregs[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_68_clk),
    .D(_00481_),
    .Q(\core.cpuregs[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_44_clk),
    .D(_00482_),
    .Q(\core.cpuregs[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_68_clk),
    .D(_00483_),
    .Q(\core.cpuregs[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_46_clk),
    .D(_00484_),
    .Q(\core.cpuregs[28][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21406_ (.CLK(clknet_leaf_43_clk),
    .D(_00485_),
    .Q(\core.cpuregs[28][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21407_ (.CLK(clknet_leaf_72_clk),
    .D(_00486_),
    .Q(\core.cpuregs[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_74_clk),
    .D(_00487_),
    .Q(\core.cpuregs[28][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21409_ (.CLK(clknet_leaf_43_clk),
    .D(_00488_),
    .Q(\core.cpuregs[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_45_clk),
    .D(_00489_),
    .Q(\core.cpuregs[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_57_clk),
    .D(_00490_),
    .Q(\core.cpuregs[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_57_clk),
    .D(_00491_),
    .Q(\core.cpuregs[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_56_clk),
    .D(_00492_),
    .Q(\core.cpuregs[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_55_clk),
    .D(_00493_),
    .Q(\core.cpuregs[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_58_clk),
    .D(_00494_),
    .Q(\core.cpuregs[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_55_clk),
    .D(_00495_),
    .Q(\core.cpuregs[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_55_clk),
    .D(_00496_),
    .Q(\core.cpuregs[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_61_clk),
    .D(_00497_),
    .Q(\core.cpuregs[28][26] ));
 sky130_fd_sc_hd__dfxtp_2 _21419_ (.CLK(clknet_leaf_62_clk),
    .D(_00498_),
    .Q(\core.cpuregs[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_57_clk),
    .D(_00499_),
    .Q(\core.cpuregs[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_69_clk),
    .D(_00500_),
    .Q(\core.cpuregs[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_61_clk),
    .D(_00501_),
    .Q(\core.cpuregs[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_70_clk),
    .D(_00502_),
    .Q(\core.cpuregs[28][31] ));
 sky130_fd_sc_hd__dfxtp_2 _21424_ (.CLK(clknet_leaf_6_clk),
    .D(_00503_),
    .Q(\core.is_alu_reg_reg ));
 sky130_fd_sc_hd__dfxtp_2 _21425_ (.CLK(clknet_leaf_18_clk),
    .D(_00504_),
    .Q(\core.is_alu_reg_imm ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_5_clk),
    .D(_00505_),
    .Q(\core.instr_auipc ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_2_clk),
    .D(_00506_),
    .Q(\core.instr_lui ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_22_clk),
    .D(\core.alu_out[0] ),
    .Q(\core.alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[1] ),
    .Q(\core.alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_0_clk),
    .D(\core.alu_out[2] ),
    .Q(\core.alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21431_ (.CLK(clknet_leaf_0_clk),
    .D(\core.alu_out[3] ),
    .Q(\core.alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_4_clk),
    .D(\core.alu_out[4] ),
    .Q(\core.alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_4 _21433_ (.CLK(clknet_leaf_4_clk),
    .D(\core.alu_out[5] ),
    .Q(\core.alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21434_ (.CLK(clknet_leaf_4_clk),
    .D(\core.alu_out[6] ),
    .Q(\core.alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(clknet_leaf_2_clk),
    .D(\core.alu_out[7] ),
    .Q(\core.alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(clknet_leaf_2_clk),
    .D(\core.alu_out[8] ),
    .Q(\core.alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[9] ),
    .Q(\core.alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(clknet_leaf_2_clk),
    .D(\core.alu_out[10] ),
    .Q(\core.alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(clknet_leaf_4_clk),
    .D(\core.alu_out[11] ),
    .Q(\core.alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(clknet_leaf_2_clk),
    .D(\core.alu_out[12] ),
    .Q(\core.alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _21441_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[13] ),
    .Q(\core.alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[14] ),
    .Q(\core.alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[15] ),
    .Q(\core.alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[16] ),
    .Q(\core.alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(clknet_leaf_0_clk),
    .D(\core.alu_out[17] ),
    .Q(\core.alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(clknet_leaf_1_clk),
    .D(\core.alu_out[18] ),
    .Q(\core.alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_4 _21447_ (.CLK(clknet_leaf_1_clk),
    .D(\core.alu_out[19] ),
    .Q(\core.alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(clknet_leaf_2_clk),
    .D(\core.alu_out[20] ),
    .Q(\core.alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(clknet_leaf_22_clk),
    .D(\core.alu_out[21] ),
    .Q(\core.alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_4 _21450_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[22] ),
    .Q(\core.alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[23] ),
    .Q(\core.alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(clknet_leaf_21_clk),
    .D(\core.alu_out[24] ),
    .Q(\core.alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(clknet_leaf_5_clk),
    .D(\core.alu_out[25] ),
    .Q(\core.alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[26] ),
    .Q(\core.alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[27] ),
    .Q(\core.alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(clknet_leaf_21_clk),
    .D(\core.alu_out[28] ),
    .Q(\core.alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[29] ),
    .Q(\core.alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(clknet_leaf_3_clk),
    .D(\core.alu_out[30] ),
    .Q(\core.alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(clknet_leaf_22_clk),
    .D(\core.alu_out[31] ),
    .Q(\core.alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(clknet_leaf_25_clk),
    .D(_00507_),
    .Q(\core.latched_is_lb ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(clknet_leaf_25_clk),
    .D(_00508_),
    .Q(\core.latched_is_lh ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(clknet_leaf_6_clk),
    .D(_00509_),
    .Q(\core.decoder_pseudo_trigger ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(clknet_leaf_22_clk),
    .D(_00510_),
    .Q(\core.latched_branch ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(clknet_leaf_21_clk),
    .D(_00511_),
    .Q(\core.latched_stalu ));
 sky130_fd_sc_hd__dfxtp_4 _21465_ (.CLK(clknet_leaf_36_clk),
    .D(_00512_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(clknet_leaf_18_clk),
    .D(_00513_),
    .Q(\core.instr_bne ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(clknet_leaf_45_clk),
    .D(_00514_),
    .Q(\core.cpuregs[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(clknet_leaf_68_clk),
    .D(_00515_),
    .Q(\core.cpuregs[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(clknet_leaf_84_clk),
    .D(_00516_),
    .Q(\core.cpuregs[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(clknet_leaf_85_clk),
    .D(_00517_),
    .Q(\core.cpuregs[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(clknet_leaf_85_clk),
    .D(_00518_),
    .Q(\core.cpuregs[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _21472_ (.CLK(clknet_leaf_67_clk),
    .D(_00519_),
    .Q(\core.cpuregs[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(clknet_leaf_85_clk),
    .D(_00520_),
    .Q(\core.cpuregs[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(clknet_leaf_74_clk),
    .D(_00521_),
    .Q(\core.cpuregs[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(clknet_leaf_71_clk),
    .D(_00522_),
    .Q(\core.cpuregs[21][8] ));
 sky130_fd_sc_hd__dfxtp_2 _21476_ (.CLK(clknet_leaf_67_clk),
    .D(_00523_),
    .Q(\core.cpuregs[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(clknet_leaf_69_clk),
    .D(_00524_),
    .Q(\core.cpuregs[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(clknet_leaf_69_clk),
    .D(_00525_),
    .Q(\core.cpuregs[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(clknet_leaf_44_clk),
    .D(_00526_),
    .Q(\core.cpuregs[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(clknet_leaf_70_clk),
    .D(_00527_),
    .Q(\core.cpuregs[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(clknet_leaf_43_clk),
    .D(_00528_),
    .Q(\core.cpuregs[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(clknet_leaf_45_clk),
    .D(_00529_),
    .Q(\core.cpuregs[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 _21483_ (.CLK(clknet_leaf_74_clk),
    .D(_00530_),
    .Q(\core.cpuregs[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(clknet_leaf_71_clk),
    .D(_00531_),
    .Q(\core.cpuregs[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(clknet_leaf_56_clk),
    .D(_00532_),
    .Q(\core.cpuregs[21][18] ));
 sky130_fd_sc_hd__dfxtp_2 _21486_ (.CLK(clknet_leaf_54_clk),
    .D(_00533_),
    .Q(\core.cpuregs[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(clknet_leaf_58_clk),
    .D(_00534_),
    .Q(\core.cpuregs[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(clknet_leaf_62_clk),
    .D(_00535_),
    .Q(\core.cpuregs[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(clknet_leaf_54_clk),
    .D(_00536_),
    .Q(\core.cpuregs[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(clknet_leaf_61_clk),
    .D(_00537_),
    .Q(\core.cpuregs[21][23] ));
 sky130_fd_sc_hd__dfxtp_2 _21491_ (.CLK(clknet_leaf_61_clk),
    .D(_00538_),
    .Q(\core.cpuregs[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(clknet_leaf_56_clk),
    .D(_00539_),
    .Q(\core.cpuregs[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(clknet_leaf_61_clk),
    .D(_00540_),
    .Q(\core.cpuregs[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(clknet_leaf_55_clk),
    .D(_00541_),
    .Q(\core.cpuregs[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(clknet_leaf_63_clk),
    .D(_00542_),
    .Q(\core.cpuregs[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(clknet_leaf_57_clk),
    .D(_00543_),
    .Q(\core.cpuregs[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_63_clk),
    .D(_00544_),
    .Q(\core.cpuregs[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_71_clk),
    .D(_00545_),
    .Q(\core.cpuregs[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_18_clk),
    .D(_00546_),
    .Q(\core.instr_jal ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_6_clk),
    .D(_00547_),
    .Q(\core.instr_beq ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_45_clk),
    .D(_00548_),
    .Q(\core.cpuregs[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 _21502_ (.CLK(clknet_leaf_69_clk),
    .D(_00549_),
    .Q(\core.cpuregs[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_82_clk),
    .D(_00550_),
    .Q(\core.cpuregs[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_84_clk),
    .D(_00551_),
    .Q(\core.cpuregs[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_84_clk),
    .D(_00552_),
    .Q(\core.cpuregs[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_82_clk),
    .D(_00553_),
    .Q(\core.cpuregs[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_82_clk),
    .D(_00554_),
    .Q(\core.cpuregs[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_82_clk),
    .D(_00555_),
    .Q(\core.cpuregs[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_67_clk),
    .D(_00556_),
    .Q(\core.cpuregs[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_67_clk),
    .D(_00557_),
    .Q(\core.cpuregs[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_68_clk),
    .D(_00558_),
    .Q(\core.cpuregs[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_46_clk),
    .D(_00559_),
    .Q(\core.cpuregs[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_72_clk),
    .D(_00560_),
    .Q(\core.cpuregs[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_44_clk),
    .D(_00561_),
    .Q(\core.cpuregs[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_73_clk),
    .D(_00562_),
    .Q(\core.cpuregs[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_73_clk),
    .D(_00563_),
    .Q(\core.cpuregs[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_74_clk),
    .D(_00564_),
    .Q(\core.cpuregs[26][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21518_ (.CLK(clknet_leaf_43_clk),
    .D(_00565_),
    .Q(\core.cpuregs[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_46_clk),
    .D(_00566_),
    .Q(\core.cpuregs[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_57_clk),
    .D(_00567_),
    .Q(\core.cpuregs[26][19] ));
 sky130_fd_sc_hd__dfxtp_2 _21521_ (.CLK(clknet_leaf_53_clk),
    .D(_00568_),
    .Q(\core.cpuregs[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_56_clk),
    .D(_00569_),
    .Q(\core.cpuregs[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_53_clk),
    .D(_00570_),
    .Q(\core.cpuregs[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_55_clk),
    .D(_00571_),
    .Q(\core.cpuregs[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_53_clk),
    .D(_00572_),
    .Q(\core.cpuregs[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_55_clk),
    .D(_00573_),
    .Q(\core.cpuregs[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_55_clk),
    .D(_00574_),
    .Q(\core.cpuregs[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_62_clk),
    .D(_00575_),
    .Q(\core.cpuregs[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_69_clk),
    .D(_00576_),
    .Q(\core.cpuregs[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_69_clk),
    .D(_00577_),
    .Q(\core.cpuregs[26][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21531_ (.CLK(clknet_leaf_69_clk),
    .D(_00578_),
    .Q(\core.cpuregs[26][30] ));
 sky130_fd_sc_hd__dfxtp_2 _21532_ (.CLK(clknet_leaf_44_clk),
    .D(_00579_),
    .Q(\core.cpuregs[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_18_clk),
    .D(_00580_),
    .Q(\core.instr_sh ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_18_clk),
    .D(_00581_),
    .Q(\core.instr_slti ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(clknet_leaf_17_clk),
    .D(_00582_),
    .Q(\core.instr_sltiu ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_18_clk),
    .D(_00583_),
    .Q(\core.instr_ori ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(clknet_leaf_21_clk),
    .D(_00584_),
    .Q(\core.latched_store ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_6_clk),
    .D(_00585_),
    .Q(\core.instr_srli ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(clknet_leaf_18_clk),
    .D(_00586_),
    .Q(\core.instr_add ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_18_clk),
    .D(_00587_),
    .Q(\core.instr_sll ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(clknet_leaf_18_clk),
    .D(_00588_),
    .Q(\core.instr_xor ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(clknet_leaf_6_clk),
    .D(_00589_),
    .Q(\core.instr_sra ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(clknet_leaf_5_clk),
    .D(_00590_),
    .Q(\core.is_compare ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_37_clk),
    .D(_00591_),
    .Q(\core.latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21545_ (.CLK(clknet_leaf_37_clk),
    .D(_00592_),
    .Q(\core.latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(clknet_leaf_37_clk),
    .D(_00593_),
    .Q(\core.latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_37_clk),
    .D(_00594_),
    .Q(\core.latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(clknet_leaf_37_clk),
    .D(_00595_),
    .Q(\core.latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_11_clk),
    .D(_00596_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(clknet_leaf_11_clk),
    .D(_00597_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_75_clk),
    .D(_00598_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(clknet_3_0__leaf_clk),
    .D(_00599_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(clknet_leaf_19_clk),
    .D(_00600_),
    .Q(\core.instr_rdcycleh ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(clknet_leaf_42_clk),
    .D(_00601_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(clknet_leaf_5_clk),
    .D(_00602_),
    .Q(\core.instr_fence ));
 sky130_fd_sc_hd__dfxtp_2 _21556_ (.CLK(clknet_leaf_20_clk),
    .D(_00603_),
    .Q(\core.mem_do_wdata ));
 sky130_fd_sc_hd__dfxtp_2 _21557_ (.CLK(clknet_leaf_18_clk),
    .D(_00030_),
    .Q(\core.decoder_trigger ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(clknet_leaf_4_clk),
    .D(_00604_),
    .Q(\core.mem_la_wdata[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21559_ (.CLK(clknet_leaf_0_clk),
    .D(_00605_),
    .Q(\core.mem_la_wdata[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(clknet_leaf_0_clk),
    .D(_00606_),
    .Q(\core.mem_la_wdata[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(clknet_leaf_0_clk),
    .D(_00607_),
    .Q(\core.mem_la_wdata[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(clknet_leaf_0_clk),
    .D(_00608_),
    .Q(\core.mem_la_wdata[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(clknet_leaf_0_clk),
    .D(_00609_),
    .Q(\core.mem_la_wdata[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(clknet_leaf_0_clk),
    .D(_00610_),
    .Q(\core.mem_la_wdata[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(clknet_leaf_0_clk),
    .D(_00611_),
    .Q(\core.mem_la_wdata[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21566_ (.CLK(clknet_leaf_79_clk),
    .D(_00612_),
    .Q(\core.pcpi_rs2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(clknet_leaf_0_clk),
    .D(_00613_),
    .Q(\core.pcpi_rs2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21568_ (.CLK(clknet_leaf_0_clk),
    .D(_00614_),
    .Q(\core.pcpi_rs2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(clknet_leaf_0_clk),
    .D(_00615_),
    .Q(\core.pcpi_rs2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(clknet_leaf_1_clk),
    .D(_00616_),
    .Q(\core.pcpi_rs2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(clknet_leaf_24_clk),
    .D(_00617_),
    .Q(\core.pcpi_rs2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _21572_ (.CLK(clknet_leaf_1_clk),
    .D(_00618_),
    .Q(\core.pcpi_rs2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(clknet_leaf_37_clk),
    .D(_00619_),
    .Q(\core.pcpi_rs2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(clknet_leaf_0_clk),
    .D(_00620_),
    .Q(\core.pcpi_rs2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(clknet_leaf_1_clk),
    .D(_00621_),
    .Q(\core.pcpi_rs2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(clknet_leaf_0_clk),
    .D(_00622_),
    .Q(\core.pcpi_rs2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _21577_ (.CLK(clknet_leaf_0_clk),
    .D(_00623_),
    .Q(\core.pcpi_rs2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21578_ (.CLK(clknet_leaf_1_clk),
    .D(_00624_),
    .Q(\core.pcpi_rs2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21579_ (.CLK(clknet_leaf_1_clk),
    .D(_00625_),
    .Q(\core.pcpi_rs2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(clknet_leaf_0_clk),
    .D(_00626_),
    .Q(\core.pcpi_rs2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _21581_ (.CLK(clknet_leaf_2_clk),
    .D(_00627_),
    .Q(\core.pcpi_rs2[23] ));
 sky130_fd_sc_hd__dfxtp_4 _21582_ (.CLK(clknet_leaf_0_clk),
    .D(_00628_),
    .Q(\core.pcpi_rs2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(clknet_leaf_1_clk),
    .D(_00629_),
    .Q(\core.pcpi_rs2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21584_ (.CLK(clknet_leaf_23_clk),
    .D(_00630_),
    .Q(\core.pcpi_rs2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21585_ (.CLK(clknet_leaf_24_clk),
    .D(_00631_),
    .Q(\core.pcpi_rs2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21586_ (.CLK(clknet_leaf_79_clk),
    .D(_00632_),
    .Q(\core.pcpi_rs2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21587_ (.CLK(clknet_leaf_24_clk),
    .D(_00633_),
    .Q(\core.pcpi_rs2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21588_ (.CLK(clknet_leaf_1_clk),
    .D(_00634_),
    .Q(\core.pcpi_rs2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21589_ (.CLK(clknet_leaf_24_clk),
    .D(_00635_),
    .Q(\core.pcpi_rs2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21590_ (.CLK(clknet_leaf_17_clk),
    .D(_00636_),
    .Q(\core.instr_bge ));
 sky130_fd_sc_hd__dfxtp_1 _21591_ (.CLK(clknet_leaf_17_clk),
    .D(_00637_),
    .Q(\core.instr_bltu ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(clknet_leaf_5_clk),
    .D(_00638_),
    .Q(\core.instr_jalr ));
 sky130_fd_sc_hd__dfxtp_2 _21593_ (.CLK(clknet_leaf_6_clk),
    .D(_00639_),
    .Q(\core.instr_lb ));
 sky130_fd_sc_hd__dfxtp_2 _21594_ (.CLK(clknet_leaf_70_clk),
    .D(_00640_),
    .Q(\core.cpuregs[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(clknet_leaf_45_clk),
    .D(_00641_),
    .Q(\core.cpuregs[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 _21596_ (.CLK(clknet_leaf_83_clk),
    .D(_00642_),
    .Q(\core.cpuregs[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21597_ (.CLK(clknet_leaf_84_clk),
    .D(_00643_),
    .Q(\core.cpuregs[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(clknet_leaf_85_clk),
    .D(_00644_),
    .Q(\core.cpuregs[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21599_ (.CLK(clknet_leaf_67_clk),
    .D(_00645_),
    .Q(\core.cpuregs[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 _21600_ (.CLK(clknet_leaf_68_clk),
    .D(_00646_),
    .Q(\core.cpuregs[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21601_ (.CLK(clknet_leaf_74_clk),
    .D(_00647_),
    .Q(\core.cpuregs[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21602_ (.CLK(clknet_leaf_70_clk),
    .D(_00648_),
    .Q(\core.cpuregs[20][8] ));
 sky130_fd_sc_hd__dfxtp_2 _21603_ (.CLK(clknet_leaf_72_clk),
    .D(_00649_),
    .Q(\core.cpuregs[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21604_ (.CLK(clknet_leaf_71_clk),
    .D(_00650_),
    .Q(\core.cpuregs[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21605_ (.CLK(clknet_leaf_70_clk),
    .D(_00651_),
    .Q(\core.cpuregs[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21606_ (.CLK(clknet_leaf_72_clk),
    .D(_00652_),
    .Q(\core.cpuregs[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_56_clk),
    .D(_00653_),
    .Q(\core.cpuregs[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_43_clk),
    .D(_00654_),
    .Q(\core.cpuregs[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21609_ (.CLK(clknet_leaf_72_clk),
    .D(_00655_),
    .Q(\core.cpuregs[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_72_clk),
    .D(_00656_),
    .Q(\core.cpuregs[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_45_clk),
    .D(_00657_),
    .Q(\core.cpuregs[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_57_clk),
    .D(_00658_),
    .Q(\core.cpuregs[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_53_clk),
    .D(_00659_),
    .Q(\core.cpuregs[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21614_ (.CLK(clknet_leaf_62_clk),
    .D(_00660_),
    .Q(\core.cpuregs[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_53_clk),
    .D(_00661_),
    .Q(\core.cpuregs[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_53_clk),
    .D(_00662_),
    .Q(\core.cpuregs[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_54_clk),
    .D(_00663_),
    .Q(\core.cpuregs[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21618_ (.CLK(clknet_leaf_54_clk),
    .D(_00664_),
    .Q(\core.cpuregs[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21619_ (.CLK(clknet_leaf_58_clk),
    .D(_00665_),
    .Q(\core.cpuregs[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_69_clk),
    .D(_00666_),
    .Q(\core.cpuregs[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_58_clk),
    .D(_00667_),
    .Q(\core.cpuregs[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_69_clk),
    .D(_00668_),
    .Q(\core.cpuregs[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_61_clk),
    .D(_00669_),
    .Q(\core.cpuregs[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_62_clk),
    .D(_00670_),
    .Q(\core.cpuregs[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_69_clk),
    .D(_00671_),
    .Q(\core.cpuregs[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21626_ (.CLK(clknet_leaf_45_clk),
    .D(_00672_),
    .Q(\core.cpuregs[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_68_clk),
    .D(_00673_),
    .Q(\core.cpuregs[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_83_clk),
    .D(_00674_),
    .Q(\core.cpuregs[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21629_ (.CLK(clknet_leaf_82_clk),
    .D(_00675_),
    .Q(\core.cpuregs[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21630_ (.CLK(clknet_leaf_85_clk),
    .D(_00676_),
    .Q(\core.cpuregs[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21631_ (.CLK(clknet_leaf_85_clk),
    .D(_00677_),
    .Q(\core.cpuregs[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21632_ (.CLK(clknet_leaf_85_clk),
    .D(_00678_),
    .Q(\core.cpuregs[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_85_clk),
    .D(_00679_),
    .Q(\core.cpuregs[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_44_clk),
    .D(_00680_),
    .Q(\core.cpuregs[25][8] ));
 sky130_fd_sc_hd__dfxtp_2 _21635_ (.CLK(clknet_leaf_74_clk),
    .D(_00681_),
    .Q(\core.cpuregs[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21636_ (.CLK(clknet_leaf_74_clk),
    .D(_00682_),
    .Q(\core.cpuregs[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_46_clk),
    .D(_00683_),
    .Q(\core.cpuregs[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21638_ (.CLK(clknet_leaf_75_clk),
    .D(_00684_),
    .Q(\core.cpuregs[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_44_clk),
    .D(_00685_),
    .Q(\core.cpuregs[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21640_ (.CLK(clknet_leaf_73_clk),
    .D(_00686_),
    .Q(\core.cpuregs[25][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21641_ (.CLK(clknet_leaf_74_clk),
    .D(_00687_),
    .Q(\core.cpuregs[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21642_ (.CLK(clknet_leaf_73_clk),
    .D(_00688_),
    .Q(\core.cpuregs[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21643_ (.CLK(clknet_leaf_42_clk),
    .D(_00689_),
    .Q(\core.cpuregs[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_46_clk),
    .D(_00690_),
    .Q(\core.cpuregs[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21645_ (.CLK(clknet_leaf_52_clk),
    .D(_00691_),
    .Q(\core.cpuregs[25][19] ));
 sky130_fd_sc_hd__dfxtp_2 _21646_ (.CLK(clknet_leaf_52_clk),
    .D(_00692_),
    .Q(\core.cpuregs[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21647_ (.CLK(clknet_leaf_55_clk),
    .D(_00693_),
    .Q(\core.cpuregs[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21648_ (.CLK(clknet_leaf_57_clk),
    .D(_00694_),
    .Q(\core.cpuregs[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21649_ (.CLK(clknet_leaf_53_clk),
    .D(_00695_),
    .Q(\core.cpuregs[25][23] ));
 sky130_fd_sc_hd__dfxtp_2 _21650_ (.CLK(clknet_leaf_71_clk),
    .D(_00696_),
    .Q(\core.cpuregs[25][24] ));
 sky130_fd_sc_hd__dfxtp_2 _21651_ (.CLK(clknet_leaf_55_clk),
    .D(_00697_),
    .Q(\core.cpuregs[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_62_clk),
    .D(_00698_),
    .Q(\core.cpuregs[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_54_clk),
    .D(_00699_),
    .Q(\core.cpuregs[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_61_clk),
    .D(_00700_),
    .Q(\core.cpuregs[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_70_clk),
    .D(_00701_),
    .Q(\core.cpuregs[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_61_clk),
    .D(_00702_),
    .Q(\core.cpuregs[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_45_clk),
    .D(_00703_),
    .Q(\core.cpuregs[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_44_clk),
    .D(_00704_),
    .Q(\core.cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_45_clk),
    .D(_00705_),
    .Q(\core.cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_82_clk),
    .D(_00706_),
    .Q(\core.cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_83_clk),
    .D(_00707_),
    .Q(\core.cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_83_clk),
    .D(_00708_),
    .Q(\core.cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_75_clk),
    .D(_00709_),
    .Q(\core.cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_75_clk),
    .D(_00710_),
    .Q(\core.cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_75_clk),
    .D(_00711_),
    .Q(\core.cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_68_clk),
    .D(_00712_),
    .Q(\core.cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _21667_ (.CLK(clknet_leaf_72_clk),
    .D(_00713_),
    .Q(\core.cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_67_clk),
    .D(_00714_),
    .Q(\core.cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_43_clk),
    .D(_00715_),
    .Q(\core.cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_72_clk),
    .D(_00716_),
    .Q(\core.cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_43_clk),
    .D(_00717_),
    .Q(\core.cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21672_ (.CLK(clknet_leaf_42_clk),
    .D(_00718_),
    .Q(\core.cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_79_clk),
    .D(_00719_),
    .Q(\core.cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _21674_ (.CLK(clknet_leaf_73_clk),
    .D(_00720_),
    .Q(\core.cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _21675_ (.CLK(clknet_leaf_47_clk),
    .D(_00721_),
    .Q(\core.cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_46_clk),
    .D(_00722_),
    .Q(\core.cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _21677_ (.CLK(clknet_leaf_50_clk),
    .D(_00723_),
    .Q(\core.cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_49_clk),
    .D(_00724_),
    .Q(\core.cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_50_clk),
    .D(_00725_),
    .Q(\core.cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_34_clk),
    .D(_00726_),
    .Q(\core.cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_49_clk),
    .D(_00727_),
    .Q(\core.cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_52_clk),
    .D(_00728_),
    .Q(\core.cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_55_clk),
    .D(_00729_),
    .Q(\core.cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_53_clk),
    .D(_00730_),
    .Q(\core.cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_44_clk),
    .D(_00731_),
    .Q(\core.cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_70_clk),
    .D(_00732_),
    .Q(\core.cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _21687_ (.CLK(clknet_leaf_70_clk),
    .D(_00733_),
    .Q(\core.cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_57_clk),
    .D(_00734_),
    .Q(\core.cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(clknet_leaf_70_clk),
    .D(_00735_),
    .Q(\core.cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(clknet_leaf_24_clk),
    .D(_00736_),
    .Q(\core.decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(clknet_leaf_37_clk),
    .D(_00737_),
    .Q(\core.decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_24_clk),
    .D(_00738_),
    .Q(\core.decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(clknet_leaf_25_clk),
    .D(_00739_),
    .Q(\core.decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(clknet_leaf_25_clk),
    .D(_00740_),
    .Q(\core.decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(clknet_leaf_23_clk),
    .D(_00741_),
    .Q(\core.decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(clknet_leaf_22_clk),
    .D(_00031_),
    .Q(\core.is_lui_auipc_jal ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_5_clk),
    .D(_00742_),
    .Q(\core.decoded_imm_j[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(clknet_leaf_5_clk),
    .D(_00743_),
    .Q(\core.decoded_imm_j[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(clknet_leaf_21_clk),
    .D(_00744_),
    .Q(\core.decoded_imm_j[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_21_clk),
    .D(_00745_),
    .Q(\core.decoded_imm_j[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_22_clk),
    .D(_00746_),
    .Q(\core.decoded_imm_j[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(clknet_leaf_21_clk),
    .D(_00747_),
    .Q(\core.decoded_imm_j[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(clknet_leaf_22_clk),
    .D(_00748_),
    .Q(\core.decoded_imm_j[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(clknet_leaf_22_clk),
    .D(_00749_),
    .Q(\core.decoded_imm_j[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21705_ (.CLK(clknet_leaf_5_clk),
    .D(_00750_),
    .Q(\core.decoded_imm_j[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(clknet_leaf_3_clk),
    .D(_00751_),
    .Q(\core.decoded_imm_j[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_18_clk),
    .D(_00752_),
    .Q(\core.decoded_imm_j[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(clknet_leaf_17_clk),
    .D(_00753_),
    .Q(\core.decoded_imm_j[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21709_ (.CLK(clknet_leaf_19_clk),
    .D(_00754_),
    .Q(\core.decoded_imm_j[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21710_ (.CLK(clknet_leaf_19_clk),
    .D(_00755_),
    .Q(\core.decoded_imm_j[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21711_ (.CLK(clknet_leaf_20_clk),
    .D(_00756_),
    .Q(\core.decoded_imm_j[15] ));
 sky130_fd_sc_hd__dfxtp_2 _21712_ (.CLK(clknet_leaf_21_clk),
    .D(_00757_),
    .Q(\core.decoded_imm_j[16] ));
 sky130_fd_sc_hd__dfxtp_2 _21713_ (.CLK(clknet_leaf_20_clk),
    .D(_00758_),
    .Q(\core.decoded_imm_j[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21714_ (.CLK(clknet_leaf_22_clk),
    .D(_00759_),
    .Q(\core.decoded_imm_j[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(clknet_leaf_20_clk),
    .D(_00760_),
    .Q(\core.decoded_imm_j[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(clknet_leaf_18_clk),
    .D(_00761_),
    .Q(\core.decoded_imm_j[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(clknet_leaf_5_clk),
    .D(_00762_),
    .Q(\core.is_lb_lh_lw_lbu_lhu ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(clknet_leaf_22_clk),
    .D(_00763_),
    .Q(\core.is_slli_srli_srai ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(clknet_leaf_22_clk),
    .D(_00764_),
    .Q(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(clknet_leaf_5_clk),
    .D(_00765_),
    .Q(\core.is_sb_sh_sw ));
 sky130_fd_sc_hd__dfxtp_1 _21721_ (.CLK(clknet_leaf_5_clk),
    .D(_00766_),
    .Q(\core.is_sll_srl_sra ));
 sky130_fd_sc_hd__dfxtp_1 _21722_ (.CLK(clknet_leaf_6_clk),
    .D(_00032_),
    .Q(\core.is_slti_blt_slt ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(clknet_leaf_17_clk),
    .D(_00033_),
    .Q(\core.is_sltiu_bltu_sltu ));
 sky130_fd_sc_hd__dfxtp_1 _21724_ (.CLK(clknet_leaf_18_clk),
    .D(_00767_),
    .Q(\core.is_beq_bne_blt_bge_bltu_bgeu ));
 sky130_fd_sc_hd__dfxtp_4 _21725_ (.CLK(clknet_leaf_23_clk),
    .D(_00768_),
    .Q(\core.decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(clknet_leaf_2_clk),
    .D(_00769_),
    .Q(\core.decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_4 _21727_ (.CLK(clknet_leaf_23_clk),
    .D(_00770_),
    .Q(\core.decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_23_clk),
    .D(_00771_),
    .Q(\core.decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_23_clk),
    .D(_00772_),
    .Q(\core.decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_22_clk),
    .D(_00773_),
    .Q(\core.decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_4 _21731_ (.CLK(clknet_leaf_24_clk),
    .D(_00774_),
    .Q(\core.decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 _21732_ (.CLK(clknet_leaf_22_clk),
    .D(_00775_),
    .Q(\core.decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(clknet_leaf_23_clk),
    .D(_00776_),
    .Q(\core.decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_4 _21734_ (.CLK(clknet_leaf_22_clk),
    .D(_00777_),
    .Q(\core.decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(clknet_leaf_24_clk),
    .D(_00778_),
    .Q(\core.decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_4 _21736_ (.CLK(clknet_leaf_24_clk),
    .D(_00779_),
    .Q(\core.decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_4 _21737_ (.CLK(clknet_leaf_22_clk),
    .D(_00780_),
    .Q(\core.decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(clknet_leaf_24_clk),
    .D(_00781_),
    .Q(\core.decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_24_clk),
    .D(_00782_),
    .Q(\core.decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(clknet_leaf_24_clk),
    .D(_00783_),
    .Q(\core.decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_4 _21741_ (.CLK(clknet_leaf_24_clk),
    .D(_00784_),
    .Q(\core.decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(clknet_leaf_22_clk),
    .D(_00785_),
    .Q(\core.decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(clknet_leaf_22_clk),
    .D(_00786_),
    .Q(\core.decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(clknet_leaf_2_clk),
    .D(_00787_),
    .Q(\core.decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21745_ (.CLK(clknet_leaf_2_clk),
    .D(_00788_),
    .Q(\core.decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(clknet_leaf_22_clk),
    .D(_00789_),
    .Q(\core.decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(clknet_leaf_2_clk),
    .D(_00790_),
    .Q(\core.decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(clknet_leaf_22_clk),
    .D(_00791_),
    .Q(\core.decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_1_clk),
    .D(_00792_),
    .Q(\core.decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_2_clk),
    .D(_00793_),
    .Q(\core.decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_2_clk),
    .D(_00794_),
    .Q(\core.decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_3_clk),
    .D(_00795_),
    .Q(\core.decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21753_ (.CLK(clknet_leaf_2_clk),
    .D(_00796_),
    .Q(\core.decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(clknet_leaf_3_clk),
    .D(_00797_),
    .Q(\core.decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(clknet_leaf_21_clk),
    .D(_00798_),
    .Q(\core.decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_44_clk),
    .D(_00799_),
    .Q(\core.cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(clknet_leaf_44_clk),
    .D(_00800_),
    .Q(\core.cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_81_clk),
    .D(_00801_),
    .Q(\core.cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(clknet_leaf_85_clk),
    .D(_00802_),
    .Q(\core.cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_83_clk),
    .D(_00803_),
    .Q(\core.cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_75_clk),
    .D(_00804_),
    .Q(\core.cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_75_clk),
    .D(_00805_),
    .Q(\core.cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_82_clk),
    .D(_00806_),
    .Q(\core.cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_71_clk),
    .D(_00807_),
    .Q(\core.cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(clknet_leaf_75_clk),
    .D(_00808_),
    .Q(\core.cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(clknet_leaf_74_clk),
    .D(_00809_),
    .Q(\core.cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21767_ (.CLK(clknet_leaf_44_clk),
    .D(_00810_),
    .Q(\core.cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(clknet_leaf_74_clk),
    .D(_00811_),
    .Q(\core.cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _21769_ (.CLK(clknet_leaf_47_clk),
    .D(_00812_),
    .Q(\core.cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(clknet_leaf_43_clk),
    .D(_00813_),
    .Q(\core.cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(clknet_leaf_42_clk),
    .D(_00814_),
    .Q(\core.cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _21772_ (.CLK(clknet_leaf_77_clk),
    .D(_00815_),
    .Q(\core.cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(clknet_leaf_42_clk),
    .D(_00816_),
    .Q(\core.cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_46_clk),
    .D(_00817_),
    .Q(\core.cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(clknet_leaf_52_clk),
    .D(_00818_),
    .Q(\core.cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _21776_ (.CLK(clknet_leaf_52_clk),
    .D(_00819_),
    .Q(\core.cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _21777_ (.CLK(clknet_leaf_57_clk),
    .D(_00820_),
    .Q(\core.cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_57_clk),
    .D(_00821_),
    .Q(\core.cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_53_clk),
    .D(_00822_),
    .Q(\core.cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_55_clk),
    .D(_00823_),
    .Q(\core.cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _21781_ (.CLK(clknet_leaf_57_clk),
    .D(_00824_),
    .Q(\core.cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _21782_ (.CLK(clknet_leaf_62_clk),
    .D(_00825_),
    .Q(\core.cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _21783_ (.CLK(clknet_leaf_62_clk),
    .D(_00826_),
    .Q(\core.cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(clknet_leaf_62_clk),
    .D(_00827_),
    .Q(\core.cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_61_clk),
    .D(_00828_),
    .Q(\core.cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21786_ (.CLK(clknet_leaf_69_clk),
    .D(_00829_),
    .Q(\core.cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(clknet_leaf_56_clk),
    .D(_00830_),
    .Q(\core.cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(clknet_leaf_42_clk),
    .D(_00831_),
    .Q(\core.cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(clknet_leaf_73_clk),
    .D(_00832_),
    .Q(\core.cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_82_clk),
    .D(_00833_),
    .Q(\core.cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(clknet_leaf_83_clk),
    .D(_00834_),
    .Q(\core.cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(clknet_leaf_83_clk),
    .D(_00835_),
    .Q(\core.cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(clknet_leaf_83_clk),
    .D(_00836_),
    .Q(\core.cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(clknet_leaf_75_clk),
    .D(_00837_),
    .Q(\core.cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(clknet_leaf_81_clk),
    .D(_00838_),
    .Q(\core.cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _21796_ (.CLK(clknet_leaf_75_clk),
    .D(_00839_),
    .Q(\core.cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_76_clk),
    .D(_00840_),
    .Q(\core.cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(clknet_leaf_76_clk),
    .D(_00841_),
    .Q(\core.cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21799_ (.CLK(clknet_leaf_73_clk),
    .D(_00842_),
    .Q(\core.cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(clknet_leaf_76_clk),
    .D(_00843_),
    .Q(\core.cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(clknet_leaf_42_clk),
    .D(_00844_),
    .Q(\core.cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(clknet_leaf_77_clk),
    .D(_00845_),
    .Q(\core.cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(clknet_leaf_42_clk),
    .D(_00846_),
    .Q(\core.cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _21804_ (.CLK(clknet_leaf_78_clk),
    .D(_00847_),
    .Q(\core.cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(clknet_leaf_39_clk),
    .D(_00848_),
    .Q(\core.cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(clknet_leaf_47_clk),
    .D(_00849_),
    .Q(\core.cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(clknet_leaf_50_clk),
    .D(_00850_),
    .Q(\core.cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(clknet_leaf_46_clk),
    .D(_00851_),
    .Q(\core.cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(clknet_leaf_50_clk),
    .D(_00852_),
    .Q(\core.cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(clknet_leaf_50_clk),
    .D(_00853_),
    .Q(\core.cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(clknet_leaf_52_clk),
    .D(_00854_),
    .Q(\core.cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(clknet_leaf_50_clk),
    .D(_00855_),
    .Q(\core.cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(clknet_leaf_52_clk),
    .D(_00856_),
    .Q(\core.cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(clknet_leaf_44_clk),
    .D(_00857_),
    .Q(\core.cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(clknet_leaf_56_clk),
    .D(_00858_),
    .Q(\core.cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _21816_ (.CLK(clknet_leaf_55_clk),
    .D(_00859_),
    .Q(\core.cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(clknet_leaf_55_clk),
    .D(_00860_),
    .Q(\core.cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(clknet_leaf_57_clk),
    .D(_00861_),
    .Q(\core.cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(clknet_leaf_47_clk),
    .D(_00862_),
    .Q(\core.cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _21820_ (.CLK(clknet_leaf_39_clk),
    .D(_00863_),
    .Q(\core.cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(clknet_leaf_73_clk),
    .D(_00864_),
    .Q(\core.cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(clknet_leaf_82_clk),
    .D(_00865_),
    .Q(\core.cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _21823_ (.CLK(clknet_leaf_83_clk),
    .D(_00866_),
    .Q(\core.cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(clknet_leaf_80_clk),
    .D(_00867_),
    .Q(\core.cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(clknet_leaf_80_clk),
    .D(_00868_),
    .Q(\core.cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(clknet_leaf_80_clk),
    .D(_00869_),
    .Q(\core.cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(clknet_leaf_79_clk),
    .D(_00870_),
    .Q(\core.cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(clknet_leaf_78_clk),
    .D(_00871_),
    .Q(\core.cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(clknet_leaf_76_clk),
    .D(_00872_),
    .Q(\core.cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(clknet_leaf_78_clk),
    .D(_00873_),
    .Q(\core.cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(clknet_leaf_37_clk),
    .D(_00874_),
    .Q(\core.cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(clknet_leaf_78_clk),
    .D(_00875_),
    .Q(\core.cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(clknet_leaf_38_clk),
    .D(_00876_),
    .Q(\core.cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(clknet_leaf_38_clk),
    .D(_00877_),
    .Q(\core.cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(clknet_leaf_40_clk),
    .D(_00878_),
    .Q(\core.cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(clknet_leaf_77_clk),
    .D(_00879_),
    .Q(\core.cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(clknet_leaf_38_clk),
    .D(_00880_),
    .Q(\core.cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(clknet_leaf_39_clk),
    .D(_00881_),
    .Q(\core.cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(clknet_leaf_41_clk),
    .D(_00882_),
    .Q(\core.cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(clknet_leaf_40_clk),
    .D(_00883_),
    .Q(\core.cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(clknet_leaf_35_clk),
    .D(_00884_),
    .Q(\core.cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(clknet_leaf_41_clk),
    .D(_00885_),
    .Q(\core.cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(clknet_leaf_35_clk),
    .D(_00886_),
    .Q(\core.cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(clknet_leaf_35_clk),
    .D(_00887_),
    .Q(\core.cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(clknet_leaf_36_clk),
    .D(_00888_),
    .Q(\core.cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _21846_ (.CLK(clknet_leaf_48_clk),
    .D(_00889_),
    .Q(\core.cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(clknet_leaf_49_clk),
    .D(_00890_),
    .Q(\core.cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _21848_ (.CLK(clknet_leaf_47_clk),
    .D(_00891_),
    .Q(\core.cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(clknet_leaf_47_clk),
    .D(_00892_),
    .Q(\core.cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(clknet_leaf_78_clk),
    .D(_00893_),
    .Q(\core.cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(clknet_leaf_42_clk),
    .D(_00894_),
    .Q(\core.cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(clknet_leaf_78_clk),
    .D(_00895_),
    .Q(\core.cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(clknet_leaf_73_clk),
    .D(_00896_),
    .Q(\core.cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(clknet_leaf_83_clk),
    .D(_00897_),
    .Q(\core.cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(clknet_leaf_80_clk),
    .D(_00898_),
    .Q(\core.cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(clknet_leaf_80_clk),
    .D(_00899_),
    .Q(\core.cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(clknet_leaf_80_clk),
    .D(_00900_),
    .Q(\core.cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(clknet_leaf_79_clk),
    .D(_00901_),
    .Q(\core.cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(clknet_leaf_80_clk),
    .D(_00902_),
    .Q(\core.cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(clknet_leaf_76_clk),
    .D(_00903_),
    .Q(\core.cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(clknet_leaf_78_clk),
    .D(_00904_),
    .Q(\core.cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(clknet_leaf_78_clk),
    .D(_00905_),
    .Q(\core.cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21863_ (.CLK(clknet_leaf_39_clk),
    .D(_00906_),
    .Q(\core.cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(clknet_leaf_78_clk),
    .D(_00907_),
    .Q(\core.cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(clknet_leaf_40_clk),
    .D(_00908_),
    .Q(\core.cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(clknet_leaf_38_clk),
    .D(_00909_),
    .Q(\core.cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(clknet_leaf_38_clk),
    .D(_00910_),
    .Q(\core.cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(clknet_leaf_38_clk),
    .D(_00911_),
    .Q(\core.cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(clknet_leaf_38_clk),
    .D(_00912_),
    .Q(\core.cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(clknet_leaf_40_clk),
    .D(_00913_),
    .Q(\core.cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(clknet_leaf_41_clk),
    .D(_00914_),
    .Q(\core.cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(clknet_leaf_40_clk),
    .D(_00915_),
    .Q(\core.cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _21873_ (.CLK(clknet_leaf_41_clk),
    .D(_00916_),
    .Q(\core.cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _21874_ (.CLK(clknet_leaf_35_clk),
    .D(_00917_),
    .Q(\core.cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(clknet_leaf_35_clk),
    .D(_00918_),
    .Q(\core.cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(clknet_leaf_40_clk),
    .D(_00919_),
    .Q(\core.cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(clknet_leaf_49_clk),
    .D(_00920_),
    .Q(\core.cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _21878_ (.CLK(clknet_leaf_42_clk),
    .D(_00921_),
    .Q(\core.cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(clknet_leaf_48_clk),
    .D(_00922_),
    .Q(\core.cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _21880_ (.CLK(clknet_leaf_47_clk),
    .D(_00923_),
    .Q(\core.cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(clknet_leaf_36_clk),
    .D(_00924_),
    .Q(\core.cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _21882_ (.CLK(clknet_leaf_48_clk),
    .D(_00925_),
    .Q(\core.cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(clknet_leaf_42_clk),
    .D(_00926_),
    .Q(\core.cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(clknet_leaf_77_clk),
    .D(_00927_),
    .Q(\core.cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(clknet_leaf_42_clk),
    .D(_00928_),
    .Q(\core.cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(clknet_leaf_82_clk),
    .D(_00929_),
    .Q(\core.cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(clknet_leaf_82_clk),
    .D(_00930_),
    .Q(\core.cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(clknet_leaf_80_clk),
    .D(_00931_),
    .Q(\core.cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(clknet_leaf_76_clk),
    .D(_00932_),
    .Q(\core.cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(clknet_leaf_80_clk),
    .D(_00933_),
    .Q(\core.cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(clknet_leaf_80_clk),
    .D(_00934_),
    .Q(\core.cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(clknet_leaf_78_clk),
    .D(_00935_),
    .Q(\core.cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(clknet_leaf_78_clk),
    .D(_00936_),
    .Q(\core.cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(clknet_leaf_77_clk),
    .D(_00937_),
    .Q(\core.cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21895_ (.CLK(clknet_leaf_38_clk),
    .D(_00938_),
    .Q(\core.cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(clknet_leaf_77_clk),
    .D(_00939_),
    .Q(\core.cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(clknet_leaf_38_clk),
    .D(_00940_),
    .Q(\core.cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21898_ (.CLK(clknet_leaf_38_clk),
    .D(_00941_),
    .Q(\core.cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(clknet_leaf_40_clk),
    .D(_00942_),
    .Q(\core.cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(clknet_leaf_38_clk),
    .D(_00943_),
    .Q(\core.cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(clknet_leaf_38_clk),
    .D(_00944_),
    .Q(\core.cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(clknet_leaf_39_clk),
    .D(_00945_),
    .Q(\core.cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(clknet_leaf_40_clk),
    .D(_00946_),
    .Q(\core.cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(clknet_leaf_40_clk),
    .D(_00947_),
    .Q(\core.cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(clknet_leaf_36_clk),
    .D(_00948_),
    .Q(\core.cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(clknet_leaf_41_clk),
    .D(_00949_),
    .Q(\core.cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(clknet_leaf_41_clk),
    .D(_00950_),
    .Q(\core.cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(clknet_leaf_40_clk),
    .D(_00951_),
    .Q(\core.cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _21909_ (.CLK(clknet_leaf_48_clk),
    .D(_00952_),
    .Q(\core.cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(clknet_leaf_41_clk),
    .D(_00953_),
    .Q(\core.cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _21911_ (.CLK(clknet_leaf_41_clk),
    .D(_00954_),
    .Q(\core.cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(clknet_leaf_48_clk),
    .D(_00955_),
    .Q(\core.cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(clknet_leaf_48_clk),
    .D(_00956_),
    .Q(\core.cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(clknet_leaf_41_clk),
    .D(_00957_),
    .Q(\core.cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _21915_ (.CLK(clknet_leaf_42_clk),
    .D(_00958_),
    .Q(\core.cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(clknet_leaf_39_clk),
    .D(_00959_),
    .Q(\core.cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(clknet_leaf_78_clk),
    .D(_00960_),
    .Q(\core.cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(clknet_leaf_83_clk),
    .D(_00961_),
    .Q(\core.cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(clknet_leaf_83_clk),
    .D(_00962_),
    .Q(\core.cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(clknet_leaf_81_clk),
    .D(_00963_),
    .Q(\core.cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(clknet_leaf_81_clk),
    .D(_00964_),
    .Q(\core.cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(clknet_leaf_80_clk),
    .D(_00965_),
    .Q(\core.cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(clknet_leaf_79_clk),
    .D(_00966_),
    .Q(\core.cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(clknet_leaf_78_clk),
    .D(_00967_),
    .Q(\core.cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(clknet_leaf_79_clk),
    .D(_00968_),
    .Q(\core.cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _21926_ (.CLK(clknet_leaf_78_clk),
    .D(_00969_),
    .Q(\core.cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(clknet_leaf_37_clk),
    .D(_00970_),
    .Q(\core.cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(clknet_leaf_78_clk),
    .D(_00971_),
    .Q(\core.cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(clknet_leaf_38_clk),
    .D(_00972_),
    .Q(\core.cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _21930_ (.CLK(clknet_leaf_38_clk),
    .D(_00973_),
    .Q(\core.cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21931_ (.CLK(clknet_leaf_38_clk),
    .D(_00974_),
    .Q(\core.cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(clknet_leaf_37_clk),
    .D(_00975_),
    .Q(\core.cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(clknet_leaf_37_clk),
    .D(_00976_),
    .Q(\core.cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(clknet_leaf_40_clk),
    .D(_00977_),
    .Q(\core.cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(clknet_leaf_40_clk),
    .D(_00978_),
    .Q(\core.cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(clknet_leaf_40_clk),
    .D(_00979_),
    .Q(\core.cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(clknet_leaf_35_clk),
    .D(_00980_),
    .Q(\core.cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(clknet_leaf_40_clk),
    .D(_00981_),
    .Q(\core.cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(clknet_leaf_35_clk),
    .D(_00982_),
    .Q(\core.cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(clknet_leaf_40_clk),
    .D(_00983_),
    .Q(\core.cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(clknet_leaf_41_clk),
    .D(_00984_),
    .Q(\core.cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(clknet_leaf_48_clk),
    .D(_00985_),
    .Q(\core.cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(clknet_leaf_41_clk),
    .D(_00986_),
    .Q(\core.cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(clknet_leaf_36_clk),
    .D(_00987_),
    .Q(\core.cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(clknet_leaf_48_clk),
    .D(_00988_),
    .Q(\core.cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(clknet_leaf_48_clk),
    .D(_00989_),
    .Q(\core.cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _21947_ (.CLK(clknet_leaf_39_clk),
    .D(_00990_),
    .Q(\core.cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(clknet_leaf_77_clk),
    .D(_00991_),
    .Q(\core.cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _21949_ (.CLK(clknet_leaf_42_clk),
    .D(_00992_),
    .Q(\core.cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(clknet_leaf_75_clk),
    .D(_00993_),
    .Q(\core.cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(clknet_leaf_81_clk),
    .D(_00994_),
    .Q(\core.cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(clknet_leaf_81_clk),
    .D(_00995_),
    .Q(\core.cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(clknet_leaf_81_clk),
    .D(_00996_),
    .Q(\core.cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(clknet_leaf_81_clk),
    .D(_00997_),
    .Q(\core.cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(clknet_leaf_81_clk),
    .D(_00998_),
    .Q(\core.cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(clknet_leaf_77_clk),
    .D(_00999_),
    .Q(\core.cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(clknet_leaf_79_clk),
    .D(_01000_),
    .Q(\core.cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _21958_ (.CLK(clknet_leaf_76_clk),
    .D(_01001_),
    .Q(\core.cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(clknet_leaf_39_clk),
    .D(_01002_),
    .Q(\core.cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _21960_ (.CLK(clknet_leaf_78_clk),
    .D(_01003_),
    .Q(\core.cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(clknet_leaf_37_clk),
    .D(_01004_),
    .Q(\core.cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(clknet_leaf_37_clk),
    .D(_01005_),
    .Q(\core.cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _21963_ (.CLK(clknet_leaf_39_clk),
    .D(_01006_),
    .Q(\core.cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(clknet_leaf_38_clk),
    .D(_01007_),
    .Q(\core.cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(clknet_leaf_37_clk),
    .D(_01008_),
    .Q(\core.cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(clknet_leaf_41_clk),
    .D(_01009_),
    .Q(\core.cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _21967_ (.CLK(clknet_leaf_35_clk),
    .D(_01010_),
    .Q(\core.cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(clknet_leaf_41_clk),
    .D(_01011_),
    .Q(\core.cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(clknet_leaf_35_clk),
    .D(_01012_),
    .Q(\core.cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(clknet_leaf_49_clk),
    .D(_01013_),
    .Q(\core.cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _21971_ (.CLK(clknet_leaf_48_clk),
    .D(_01014_),
    .Q(\core.cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(clknet_leaf_41_clk),
    .D(_01015_),
    .Q(\core.cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(clknet_leaf_49_clk),
    .D(_01016_),
    .Q(\core.cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(clknet_leaf_36_clk),
    .D(_01017_),
    .Q(\core.cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(clknet_leaf_49_clk),
    .D(_01018_),
    .Q(\core.cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(clknet_leaf_50_clk),
    .D(_01019_),
    .Q(\core.cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(clknet_leaf_48_clk),
    .D(_01020_),
    .Q(\core.cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(clknet_leaf_48_clk),
    .D(_01021_),
    .Q(\core.cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(clknet_leaf_47_clk),
    .D(_01022_),
    .Q(\core.cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(clknet_leaf_77_clk),
    .D(_01023_),
    .Q(\core.cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(clknet_leaf_73_clk),
    .D(_01024_),
    .Q(\core.cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(clknet_leaf_75_clk),
    .D(_01025_),
    .Q(\core.cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(clknet_leaf_82_clk),
    .D(_01026_),
    .Q(\core.cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(clknet_leaf_81_clk),
    .D(_01027_),
    .Q(\core.cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(clknet_leaf_81_clk),
    .D(_01028_),
    .Q(\core.cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(clknet_leaf_79_clk),
    .D(_01029_),
    .Q(\core.cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(clknet_leaf_80_clk),
    .D(_01030_),
    .Q(\core.cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(clknet_leaf_76_clk),
    .D(_01031_),
    .Q(\core.cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(clknet_leaf_76_clk),
    .D(_01032_),
    .Q(\core.cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(clknet_leaf_76_clk),
    .D(_01033_),
    .Q(\core.cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _21991_ (.CLK(clknet_leaf_39_clk),
    .D(_01034_),
    .Q(\core.cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _21992_ (.CLK(clknet_leaf_78_clk),
    .D(_01035_),
    .Q(\core.cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(clknet_leaf_39_clk),
    .D(_01036_),
    .Q(\core.cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(clknet_leaf_40_clk),
    .D(_01037_),
    .Q(\core.cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(clknet_leaf_39_clk),
    .D(_01038_),
    .Q(\core.cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(clknet_leaf_38_clk),
    .D(_01039_),
    .Q(\core.cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(clknet_leaf_38_clk),
    .D(_01040_),
    .Q(\core.cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _21998_ (.CLK(clknet_leaf_40_clk),
    .D(_01041_),
    .Q(\core.cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(clknet_leaf_35_clk),
    .D(_01042_),
    .Q(\core.cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(clknet_leaf_41_clk),
    .D(_01043_),
    .Q(\core.cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(clknet_leaf_35_clk),
    .D(_01044_),
    .Q(\core.cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(clknet_leaf_36_clk),
    .D(_01045_),
    .Q(\core.cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(clknet_leaf_48_clk),
    .D(_01046_),
    .Q(\core.cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(clknet_leaf_35_clk),
    .D(_01047_),
    .Q(\core.cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(clknet_leaf_35_clk),
    .D(_01048_),
    .Q(\core.cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(clknet_leaf_36_clk),
    .D(_01049_),
    .Q(\core.cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(clknet_leaf_36_clk),
    .D(_01050_),
    .Q(\core.cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(clknet_leaf_47_clk),
    .D(_01051_),
    .Q(\core.cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(clknet_leaf_50_clk),
    .D(_01052_),
    .Q(\core.cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(clknet_leaf_36_clk),
    .D(_01053_),
    .Q(\core.cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(clknet_leaf_48_clk),
    .D(_01054_),
    .Q(\core.cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _22012_ (.CLK(clknet_leaf_73_clk),
    .D(_01055_),
    .Q(\core.cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22013_ (.CLK(clknet_leaf_43_clk),
    .D(_01056_),
    .Q(\core.cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(clknet_leaf_83_clk),
    .D(_01057_),
    .Q(\core.cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(clknet_leaf_82_clk),
    .D(_01058_),
    .Q(\core.cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(clknet_leaf_81_clk),
    .D(_01059_),
    .Q(\core.cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(clknet_leaf_75_clk),
    .D(_01060_),
    .Q(\core.cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(clknet_leaf_76_clk),
    .D(_01061_),
    .Q(\core.cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(clknet_leaf_75_clk),
    .D(_01062_),
    .Q(\core.cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(clknet_leaf_68_clk),
    .D(_01063_),
    .Q(\core.cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(clknet_leaf_68_clk),
    .D(_01064_),
    .Q(\core.cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _22022_ (.CLK(clknet_leaf_71_clk),
    .D(_01065_),
    .Q(\core.cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(clknet_leaf_43_clk),
    .D(_01066_),
    .Q(\core.cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(clknet_leaf_72_clk),
    .D(_01067_),
    .Q(\core.cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(clknet_leaf_42_clk),
    .D(_01068_),
    .Q(\core.cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(clknet_leaf_78_clk),
    .D(_01069_),
    .Q(\core.cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(clknet_leaf_47_clk),
    .D(_01070_),
    .Q(\core.cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(clknet_leaf_73_clk),
    .D(_01071_),
    .Q(\core.cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(clknet_leaf_47_clk),
    .D(_01072_),
    .Q(\core.cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(clknet_leaf_47_clk),
    .D(_01073_),
    .Q(\core.cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(clknet_leaf_50_clk),
    .D(_01074_),
    .Q(\core.cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(clknet_leaf_49_clk),
    .D(_01075_),
    .Q(\core.cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(clknet_leaf_52_clk),
    .D(_01076_),
    .Q(\core.cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(clknet_leaf_49_clk),
    .D(_01077_),
    .Q(\core.cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(clknet_leaf_50_clk),
    .D(_01078_),
    .Q(\core.cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(clknet_leaf_51_clk),
    .D(_01079_),
    .Q(\core.cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(clknet_leaf_49_clk),
    .D(_01080_),
    .Q(\core.cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(clknet_leaf_61_clk),
    .D(_01081_),
    .Q(\core.cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(clknet_leaf_52_clk),
    .D(_01082_),
    .Q(\core.cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(clknet_leaf_57_clk),
    .D(_01083_),
    .Q(\core.cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(clknet_leaf_56_clk),
    .D(_01084_),
    .Q(\core.cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(clknet_leaf_53_clk),
    .D(_01085_),
    .Q(\core.cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(clknet_leaf_70_clk),
    .D(_01086_),
    .Q(\core.cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(clknet_leaf_39_clk),
    .D(_01087_),
    .Q(\core.cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(clknet_leaf_43_clk),
    .D(_01088_),
    .Q(\core.cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(clknet_leaf_83_clk),
    .D(_01089_),
    .Q(\core.cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(clknet_leaf_83_clk),
    .D(_01090_),
    .Q(\core.cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(clknet_leaf_83_clk),
    .D(_01091_),
    .Q(\core.cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(clknet_leaf_81_clk),
    .D(_01092_),
    .Q(\core.cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(clknet_leaf_80_clk),
    .D(_01093_),
    .Q(\core.cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(clknet_leaf_80_clk),
    .D(_01094_),
    .Q(\core.cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22052_ (.CLK(clknet_leaf_76_clk),
    .D(_01095_),
    .Q(\core.cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(clknet_leaf_76_clk),
    .D(_01096_),
    .Q(\core.cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(clknet_leaf_76_clk),
    .D(_01097_),
    .Q(\core.cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22055_ (.CLK(clknet_leaf_37_clk),
    .D(_01098_),
    .Q(\core.cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(clknet_leaf_78_clk),
    .D(_01099_),
    .Q(\core.cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(clknet_leaf_40_clk),
    .D(_01100_),
    .Q(\core.cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _22058_ (.CLK(clknet_leaf_38_clk),
    .D(_01101_),
    .Q(\core.cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(clknet_leaf_39_clk),
    .D(_01102_),
    .Q(\core.cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(clknet_leaf_38_clk),
    .D(_01103_),
    .Q(\core.cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(clknet_leaf_38_clk),
    .D(_01104_),
    .Q(\core.cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(clknet_leaf_40_clk),
    .D(_01105_),
    .Q(\core.cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(clknet_leaf_35_clk),
    .D(_01106_),
    .Q(\core.cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(clknet_leaf_41_clk),
    .D(_01107_),
    .Q(\core.cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(clknet_leaf_48_clk),
    .D(_01108_),
    .Q(\core.cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(clknet_leaf_40_clk),
    .D(_01109_),
    .Q(\core.cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(clknet_leaf_48_clk),
    .D(_01110_),
    .Q(\core.cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _22068_ (.CLK(clknet_leaf_35_clk),
    .D(_01111_),
    .Q(\core.cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(clknet_leaf_49_clk),
    .D(_01112_),
    .Q(\core.cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(clknet_leaf_47_clk),
    .D(_01113_),
    .Q(\core.cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(clknet_leaf_41_clk),
    .D(_01114_),
    .Q(\core.cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(clknet_leaf_47_clk),
    .D(_01115_),
    .Q(\core.cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(clknet_leaf_49_clk),
    .D(_01116_),
    .Q(\core.cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22074_ (.CLK(clknet_leaf_48_clk),
    .D(_01117_),
    .Q(\core.cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22075_ (.CLK(clknet_leaf_42_clk),
    .D(_01118_),
    .Q(\core.cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _22076_ (.CLK(clknet_leaf_76_clk),
    .D(_01119_),
    .Q(\core.cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22077_ (.CLK(clknet_leaf_77_clk),
    .D(_01120_),
    .Q(\core.cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22078_ (.CLK(clknet_leaf_81_clk),
    .D(_01121_),
    .Q(\core.cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22079_ (.CLK(clknet_leaf_81_clk),
    .D(_01122_),
    .Q(\core.cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22080_ (.CLK(clknet_leaf_81_clk),
    .D(_01123_),
    .Q(\core.cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22081_ (.CLK(clknet_leaf_76_clk),
    .D(_01124_),
    .Q(\core.cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22082_ (.CLK(clknet_leaf_76_clk),
    .D(_01125_),
    .Q(\core.cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22083_ (.CLK(clknet_leaf_80_clk),
    .D(_01126_),
    .Q(\core.cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22084_ (.CLK(clknet_leaf_77_clk),
    .D(_01127_),
    .Q(\core.cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _22085_ (.CLK(clknet_leaf_76_clk),
    .D(_01128_),
    .Q(\core.cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22086_ (.CLK(clknet_leaf_76_clk),
    .D(_01129_),
    .Q(\core.cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22087_ (.CLK(clknet_leaf_39_clk),
    .D(_01130_),
    .Q(\core.cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22088_ (.CLK(clknet_leaf_77_clk),
    .D(_01131_),
    .Q(\core.cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22089_ (.CLK(clknet_leaf_39_clk),
    .D(_01132_),
    .Q(\core.cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _22090_ (.CLK(clknet_leaf_39_clk),
    .D(_01133_),
    .Q(\core.cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22091_ (.CLK(clknet_leaf_39_clk),
    .D(_01134_),
    .Q(\core.cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _22092_ (.CLK(clknet_leaf_77_clk),
    .D(_01135_),
    .Q(\core.cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22093_ (.CLK(clknet_leaf_41_clk),
    .D(_01136_),
    .Q(\core.cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _22094_ (.CLK(clknet_leaf_41_clk),
    .D(_01137_),
    .Q(\core.cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22095_ (.CLK(clknet_leaf_47_clk),
    .D(_01138_),
    .Q(\core.cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22096_ (.CLK(clknet_leaf_50_clk),
    .D(_01139_),
    .Q(\core.cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _22097_ (.CLK(clknet_leaf_49_clk),
    .D(_01140_),
    .Q(\core.cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _22098_ (.CLK(clknet_leaf_47_clk),
    .D(_01141_),
    .Q(\core.cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22099_ (.CLK(clknet_leaf_35_clk),
    .D(_01142_),
    .Q(\core.cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22100_ (.CLK(clknet_leaf_35_clk),
    .D(_01143_),
    .Q(\core.cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22101_ (.CLK(clknet_leaf_35_clk),
    .D(_01144_),
    .Q(\core.cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22102_ (.CLK(clknet_leaf_79_clk),
    .D(_01145_),
    .Q(\core.cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22103_ (.CLK(clknet_leaf_50_clk),
    .D(_01146_),
    .Q(\core.cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _22104_ (.CLK(clknet_leaf_46_clk),
    .D(_01147_),
    .Q(\core.cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _22105_ (.CLK(clknet_leaf_47_clk),
    .D(_01148_),
    .Q(\core.cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22106_ (.CLK(clknet_leaf_50_clk),
    .D(_01149_),
    .Q(\core.cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _22107_ (.CLK(clknet_leaf_47_clk),
    .D(_01150_),
    .Q(\core.cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22108_ (.CLK(clknet_leaf_73_clk),
    .D(_01151_),
    .Q(\core.cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22109_ (.CLK(clknet_leaf_77_clk),
    .D(_01152_),
    .Q(\core.cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22110_ (.CLK(clknet_leaf_80_clk),
    .D(_01153_),
    .Q(\core.cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22111_ (.CLK(clknet_leaf_83_clk),
    .D(_01154_),
    .Q(\core.cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22112_ (.CLK(clknet_leaf_80_clk),
    .D(_01155_),
    .Q(\core.cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22113_ (.CLK(clknet_leaf_76_clk),
    .D(_01156_),
    .Q(\core.cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22114_ (.CLK(clknet_leaf_81_clk),
    .D(_01157_),
    .Q(\core.cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22115_ (.CLK(clknet_leaf_80_clk),
    .D(_01158_),
    .Q(\core.cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22116_ (.CLK(clknet_leaf_77_clk),
    .D(_01159_),
    .Q(\core.cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _22117_ (.CLK(clknet_leaf_81_clk),
    .D(_01160_),
    .Q(\core.cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _22118_ (.CLK(clknet_leaf_76_clk),
    .D(_01161_),
    .Q(\core.cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22119_ (.CLK(clknet_leaf_39_clk),
    .D(_01162_),
    .Q(\core.cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22120_ (.CLK(clknet_leaf_76_clk),
    .D(_01163_),
    .Q(\core.cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22121_ (.CLK(clknet_leaf_39_clk),
    .D(_01164_),
    .Q(\core.cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22122_ (.CLK(clknet_leaf_38_clk),
    .D(_01165_),
    .Q(\core.cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22123_ (.CLK(clknet_leaf_39_clk),
    .D(_01166_),
    .Q(\core.cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22124_ (.CLK(clknet_leaf_38_clk),
    .D(_01167_),
    .Q(\core.cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22125_ (.CLK(clknet_leaf_40_clk),
    .D(_01168_),
    .Q(\core.cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22126_ (.CLK(clknet_leaf_41_clk),
    .D(_01169_),
    .Q(\core.cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22127_ (.CLK(clknet_leaf_48_clk),
    .D(_01170_),
    .Q(\core.cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22128_ (.CLK(clknet_leaf_49_clk),
    .D(_01171_),
    .Q(\core.cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _22129_ (.CLK(clknet_leaf_35_clk),
    .D(_01172_),
    .Q(\core.cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _22130_ (.CLK(clknet_leaf_35_clk),
    .D(_01173_),
    .Q(\core.cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22131_ (.CLK(clknet_leaf_49_clk),
    .D(_01174_),
    .Q(\core.cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22132_ (.CLK(clknet_leaf_49_clk),
    .D(_01175_),
    .Q(\core.cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22133_ (.CLK(clknet_leaf_50_clk),
    .D(_01176_),
    .Q(\core.cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22134_ (.CLK(clknet_leaf_46_clk),
    .D(_01177_),
    .Q(\core.cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _22135_ (.CLK(clknet_leaf_50_clk),
    .D(_01178_),
    .Q(\core.cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _22136_ (.CLK(clknet_leaf_50_clk),
    .D(_01179_),
    .Q(\core.cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _22137_ (.CLK(clknet_leaf_50_clk),
    .D(_01180_),
    .Q(\core.cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22138_ (.CLK(clknet_leaf_79_clk),
    .D(_01181_),
    .Q(\core.cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _22139_ (.CLK(clknet_leaf_47_clk),
    .D(_01182_),
    .Q(\core.cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22140_ (.CLK(clknet_leaf_77_clk),
    .D(_01183_),
    .Q(\core.cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22141_ (.CLK(clknet_leaf_42_clk),
    .D(_01184_),
    .Q(\core.cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22142_ (.CLK(clknet_leaf_81_clk),
    .D(_01185_),
    .Q(\core.cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22143_ (.CLK(clknet_leaf_82_clk),
    .D(_01186_),
    .Q(\core.cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _22144_ (.CLK(clknet_leaf_80_clk),
    .D(_01187_),
    .Q(\core.cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22145_ (.CLK(clknet_leaf_75_clk),
    .D(_01188_),
    .Q(\core.cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22146_ (.CLK(clknet_leaf_81_clk),
    .D(_01189_),
    .Q(\core.cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22147_ (.CLK(clknet_leaf_81_clk),
    .D(_01190_),
    .Q(\core.cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22148_ (.CLK(clknet_leaf_77_clk),
    .D(_01191_),
    .Q(\core.cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22149_ (.CLK(clknet_leaf_80_clk),
    .D(_01192_),
    .Q(\core.cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22150_ (.CLK(clknet_leaf_77_clk),
    .D(_01193_),
    .Q(\core.cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22151_ (.CLK(clknet_leaf_42_clk),
    .D(_01194_),
    .Q(\core.cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22152_ (.CLK(clknet_leaf_77_clk),
    .D(_01195_),
    .Q(\core.cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _22153_ (.CLK(clknet_leaf_42_clk),
    .D(_01196_),
    .Q(\core.cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22154_ (.CLK(clknet_leaf_40_clk),
    .D(_01197_),
    .Q(\core.cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22155_ (.CLK(clknet_leaf_43_clk),
    .D(_01198_),
    .Q(\core.cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22156_ (.CLK(clknet_leaf_77_clk),
    .D(_01199_),
    .Q(\core.cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22157_ (.CLK(clknet_leaf_39_clk),
    .D(_01200_),
    .Q(\core.cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22158_ (.CLK(clknet_leaf_42_clk),
    .D(_01201_),
    .Q(\core.cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22159_ (.CLK(clknet_leaf_49_clk),
    .D(_01202_),
    .Q(\core.cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22160_ (.CLK(clknet_leaf_49_clk),
    .D(_01203_),
    .Q(\core.cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22161_ (.CLK(clknet_leaf_49_clk),
    .D(_01204_),
    .Q(\core.cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22162_ (.CLK(clknet_leaf_34_clk),
    .D(_01205_),
    .Q(\core.cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22163_ (.CLK(clknet_leaf_49_clk),
    .D(_01206_),
    .Q(\core.cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _22164_ (.CLK(clknet_leaf_50_clk),
    .D(_01207_),
    .Q(\core.cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22165_ (.CLK(clknet_leaf_35_clk),
    .D(_01208_),
    .Q(\core.cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22166_ (.CLK(clknet_leaf_50_clk),
    .D(_01209_),
    .Q(\core.cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22167_ (.CLK(clknet_leaf_49_clk),
    .D(_01210_),
    .Q(\core.cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22168_ (.CLK(clknet_leaf_79_clk),
    .D(_01211_),
    .Q(\core.cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _22169_ (.CLK(clknet_leaf_50_clk),
    .D(_01212_),
    .Q(\core.cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22170_ (.CLK(clknet_leaf_50_clk),
    .D(_01213_),
    .Q(\core.cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22171_ (.CLK(clknet_leaf_43_clk),
    .D(_01214_),
    .Q(\core.cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22172_ (.CLK(clknet_leaf_73_clk),
    .D(_01215_),
    .Q(\core.cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22173_ (.CLK(clknet_leaf_73_clk),
    .D(_01216_),
    .Q(\core.cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22174_ (.CLK(clknet_leaf_81_clk),
    .D(_01217_),
    .Q(\core.cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22175_ (.CLK(clknet_leaf_82_clk),
    .D(_01218_),
    .Q(\core.cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _22176_ (.CLK(clknet_leaf_83_clk),
    .D(_01219_),
    .Q(\core.cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22177_ (.CLK(clknet_leaf_75_clk),
    .D(_01220_),
    .Q(\core.cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22178_ (.CLK(clknet_leaf_81_clk),
    .D(_01221_),
    .Q(\core.cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22179_ (.CLK(clknet_leaf_80_clk),
    .D(_01222_),
    .Q(\core.cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22180_ (.CLK(clknet_leaf_77_clk),
    .D(_01223_),
    .Q(\core.cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _22181_ (.CLK(clknet_leaf_76_clk),
    .D(_01224_),
    .Q(\core.cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22182_ (.CLK(clknet_leaf_77_clk),
    .D(_01225_),
    .Q(\core.cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22183_ (.CLK(clknet_leaf_78_clk),
    .D(_01226_),
    .Q(\core.cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22184_ (.CLK(clknet_leaf_77_clk),
    .D(_01227_),
    .Q(\core.cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _22185_ (.CLK(clknet_leaf_41_clk),
    .D(_01228_),
    .Q(\core.cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22186_ (.CLK(clknet_leaf_39_clk),
    .D(_01229_),
    .Q(\core.cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _22187_ (.CLK(clknet_leaf_42_clk),
    .D(_01230_),
    .Q(\core.cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22188_ (.CLK(clknet_leaf_77_clk),
    .D(_01231_),
    .Q(\core.cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _22189_ (.CLK(clknet_leaf_39_clk),
    .D(_01232_),
    .Q(\core.cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22190_ (.CLK(clknet_leaf_42_clk),
    .D(_01233_),
    .Q(\core.cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22191_ (.CLK(clknet_leaf_49_clk),
    .D(_01234_),
    .Q(\core.cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22192_ (.CLK(clknet_leaf_49_clk),
    .D(_01235_),
    .Q(\core.cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22193_ (.CLK(clknet_leaf_51_clk),
    .D(_01236_),
    .Q(\core.cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22194_ (.CLK(clknet_leaf_35_clk),
    .D(_01237_),
    .Q(\core.cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22195_ (.CLK(clknet_leaf_34_clk),
    .D(_01238_),
    .Q(\core.cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22196_ (.CLK(clknet_leaf_35_clk),
    .D(_01239_),
    .Q(\core.cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _22197_ (.CLK(clknet_leaf_50_clk),
    .D(_01240_),
    .Q(\core.cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22198_ (.CLK(clknet_leaf_46_clk),
    .D(_01241_),
    .Q(\core.cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22199_ (.CLK(clknet_leaf_34_clk),
    .D(_01242_),
    .Q(\core.cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22200_ (.CLK(clknet_leaf_50_clk),
    .D(_01243_),
    .Q(\core.cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _22201_ (.CLK(clknet_leaf_50_clk),
    .D(_01244_),
    .Q(\core.cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22202_ (.CLK(clknet_leaf_50_clk),
    .D(_01245_),
    .Q(\core.cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22203_ (.CLK(clknet_leaf_47_clk),
    .D(_01246_),
    .Q(\core.cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22204_ (.CLK(clknet_leaf_21_clk),
    .D(_00017_),
    .Q(\core.mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22205_ (.CLK(clknet_leaf_21_clk),
    .D(_00018_),
    .Q(\core.mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22206_ (.CLK(clknet_leaf_21_clk),
    .D(_00019_),
    .Q(\core.mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22207_ (.CLK(clknet_leaf_71_clk),
    .D(_01247_),
    .Q(\core.cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22208_ (.CLK(clknet_leaf_46_clk),
    .D(_01248_),
    .Q(\core.cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22209_ (.CLK(clknet_leaf_85_clk),
    .D(_01249_),
    .Q(\core.cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22210_ (.CLK(clknet_leaf_84_clk),
    .D(_01250_),
    .Q(\core.cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22211_ (.CLK(clknet_leaf_83_clk),
    .D(_01251_),
    .Q(\core.cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22212_ (.CLK(clknet_leaf_75_clk),
    .D(_01252_),
    .Q(\core.cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22213_ (.CLK(clknet_leaf_75_clk),
    .D(_01253_),
    .Q(\core.cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22214_ (.CLK(clknet_leaf_75_clk),
    .D(_01254_),
    .Q(\core.cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22215_ (.CLK(clknet_leaf_68_clk),
    .D(_01255_),
    .Q(\core.cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22216_ (.CLK(clknet_leaf_74_clk),
    .D(_01256_),
    .Q(\core.cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22217_ (.CLK(clknet_leaf_71_clk),
    .D(_01257_),
    .Q(\core.cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22218_ (.CLK(clknet_leaf_47_clk),
    .D(_01258_),
    .Q(\core.cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22219_ (.CLK(clknet_leaf_68_clk),
    .D(_01259_),
    .Q(\core.cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _22220_ (.CLK(clknet_leaf_47_clk),
    .D(_01260_),
    .Q(\core.cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22221_ (.CLK(clknet_leaf_43_clk),
    .D(_01261_),
    .Q(\core.cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22222_ (.CLK(clknet_leaf_47_clk),
    .D(_01262_),
    .Q(\core.cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22223_ (.CLK(clknet_leaf_73_clk),
    .D(_01263_),
    .Q(\core.cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22224_ (.CLK(clknet_leaf_42_clk),
    .D(_01264_),
    .Q(\core.cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _22225_ (.CLK(clknet_leaf_46_clk),
    .D(_01265_),
    .Q(\core.cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22226_ (.CLK(clknet_leaf_52_clk),
    .D(_01266_),
    .Q(\core.cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22227_ (.CLK(clknet_leaf_49_clk),
    .D(_01267_),
    .Q(\core.cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22228_ (.CLK(clknet_leaf_52_clk),
    .D(_01268_),
    .Q(\core.cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22229_ (.CLK(clknet_leaf_34_clk),
    .D(_01269_),
    .Q(\core.cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22230_ (.CLK(clknet_leaf_49_clk),
    .D(_01270_),
    .Q(\core.cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_4 _22231_ (.CLK(clknet_leaf_52_clk),
    .D(_01271_),
    .Q(\core.cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22232_ (.CLK(clknet_leaf_61_clk),
    .D(_01272_),
    .Q(\core.cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22233_ (.CLK(clknet_leaf_61_clk),
    .D(_01273_),
    .Q(\core.cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22234_ (.CLK(clknet_leaf_57_clk),
    .D(_01274_),
    .Q(\core.cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22235_ (.CLK(clknet_leaf_70_clk),
    .D(_01275_),
    .Q(\core.cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22236_ (.CLK(clknet_leaf_53_clk),
    .D(_01276_),
    .Q(\core.cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22237_ (.CLK(clknet_leaf_61_clk),
    .D(_01277_),
    .Q(\core.cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22238_ (.CLK(clknet_leaf_45_clk),
    .D(_01278_),
    .Q(\core.cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22239_ (.CLK(clknet_leaf_19_clk),
    .D(_00010_),
    .Q(\core.cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22240_ (.CLK(clknet_leaf_6_clk),
    .D(_00011_),
    .Q(\core.cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22241_ (.CLK(clknet_leaf_21_clk),
    .D(_00012_),
    .Q(\core.cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22242_ (.CLK(clknet_leaf_21_clk),
    .D(_00013_),
    .Q(\core.cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22243_ (.CLK(clknet_leaf_3_clk),
    .D(_00014_),
    .Q(\core.cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22244_ (.CLK(clknet_leaf_18_clk),
    .D(_00015_),
    .Q(\core.cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22245_ (.CLK(clknet_leaf_21_clk),
    .D(_00016_),
    .Q(\core.cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22246_ (.CLK(clknet_leaf_46_clk),
    .D(_01279_),
    .Q(\core.cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22247_ (.CLK(clknet_leaf_72_clk),
    .D(_01280_),
    .Q(\core.cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22248_ (.CLK(clknet_leaf_85_clk),
    .D(_01281_),
    .Q(\core.cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22249_ (.CLK(clknet_leaf_85_clk),
    .D(_01282_),
    .Q(\core.cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22250_ (.CLK(clknet_leaf_83_clk),
    .D(_01283_),
    .Q(\core.cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22251_ (.CLK(clknet_leaf_67_clk),
    .D(_01284_),
    .Q(\core.cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22252_ (.CLK(clknet_leaf_67_clk),
    .D(_01285_),
    .Q(\core.cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22253_ (.CLK(clknet_leaf_81_clk),
    .D(_01286_),
    .Q(\core.cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22254_ (.CLK(clknet_leaf_71_clk),
    .D(_01287_),
    .Q(\core.cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22255_ (.CLK(clknet_leaf_72_clk),
    .D(_01288_),
    .Q(\core.cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22256_ (.CLK(clknet_leaf_68_clk),
    .D(_01289_),
    .Q(\core.cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22257_ (.CLK(clknet_leaf_45_clk),
    .D(_01290_),
    .Q(\core.cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22258_ (.CLK(clknet_leaf_44_clk),
    .D(_01291_),
    .Q(\core.cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22259_ (.CLK(clknet_leaf_46_clk),
    .D(_01292_),
    .Q(\core.cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22260_ (.CLK(clknet_leaf_42_clk),
    .D(_01293_),
    .Q(\core.cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_4 _22261_ (.CLK(clknet_leaf_73_clk),
    .D(_01294_),
    .Q(\core.cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22262_ (.CLK(clknet_leaf_73_clk),
    .D(_01295_),
    .Q(\core.cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22263_ (.CLK(clknet_leaf_43_clk),
    .D(_01296_),
    .Q(\core.cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _22264_ (.CLK(clknet_leaf_55_clk),
    .D(_01297_),
    .Q(\core.cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22265_ (.CLK(clknet_leaf_52_clk),
    .D(_01298_),
    .Q(\core.cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _22266_ (.CLK(clknet_leaf_56_clk),
    .D(_01299_),
    .Q(\core.cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22267_ (.CLK(clknet_leaf_61_clk),
    .D(_01300_),
    .Q(\core.cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22268_ (.CLK(clknet_leaf_52_clk),
    .D(_01301_),
    .Q(\core.cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _22269_ (.CLK(clknet_leaf_53_clk),
    .D(_01302_),
    .Q(\core.cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22270_ (.CLK(clknet_leaf_70_clk),
    .D(_01303_),
    .Q(\core.cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22271_ (.CLK(clknet_leaf_61_clk),
    .D(_01304_),
    .Q(\core.cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22272_ (.CLK(clknet_leaf_62_clk),
    .D(_01305_),
    .Q(\core.cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22273_ (.CLK(clknet_leaf_54_clk),
    .D(_01306_),
    .Q(\core.cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22274_ (.CLK(clknet_leaf_69_clk),
    .D(_01307_),
    .Q(\core.cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22275_ (.CLK(clknet_leaf_55_clk),
    .D(_01308_),
    .Q(\core.cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _22276_ (.CLK(clknet_leaf_61_clk),
    .D(_01309_),
    .Q(\core.cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _22277_ (.CLK(clknet_leaf_71_clk),
    .D(_01310_),
    .Q(\core.cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22278_ (.CLK(clknet_leaf_45_clk),
    .D(_01311_),
    .Q(\core.cpuregs[31][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22279_ (.CLK(clknet_leaf_56_clk),
    .D(_01312_),
    .Q(\core.cpuregs[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22280_ (.CLK(clknet_leaf_82_clk),
    .D(_01313_),
    .Q(\core.cpuregs[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22281_ (.CLK(clknet_leaf_85_clk),
    .D(_01314_),
    .Q(\core.cpuregs[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22282_ (.CLK(clknet_leaf_82_clk),
    .D(_01315_),
    .Q(\core.cpuregs[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22283_ (.CLK(clknet_leaf_74_clk),
    .D(_01316_),
    .Q(\core.cpuregs[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22284_ (.CLK(clknet_leaf_74_clk),
    .D(_01317_),
    .Q(\core.cpuregs[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22285_ (.CLK(clknet_leaf_67_clk),
    .D(_01318_),
    .Q(\core.cpuregs[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22286_ (.CLK(clknet_leaf_70_clk),
    .D(_01319_),
    .Q(\core.cpuregs[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22287_ (.CLK(clknet_leaf_68_clk),
    .D(_01320_),
    .Q(\core.cpuregs[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22288_ (.CLK(clknet_leaf_68_clk),
    .D(_01321_),
    .Q(\core.cpuregs[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22289_ (.CLK(clknet_leaf_71_clk),
    .D(_01322_),
    .Q(\core.cpuregs[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22290_ (.CLK(clknet_leaf_71_clk),
    .D(_01323_),
    .Q(\core.cpuregs[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22291_ (.CLK(clknet_leaf_45_clk),
    .D(_01324_),
    .Q(\core.cpuregs[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22292_ (.CLK(clknet_leaf_72_clk),
    .D(_01325_),
    .Q(\core.cpuregs[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 _22293_ (.CLK(clknet_leaf_43_clk),
    .D(_01326_),
    .Q(\core.cpuregs[31][15] ));
 sky130_fd_sc_hd__dfxtp_2 _22294_ (.CLK(clknet_leaf_72_clk),
    .D(_01327_),
    .Q(\core.cpuregs[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22295_ (.CLK(clknet_leaf_43_clk),
    .D(_01328_),
    .Q(\core.cpuregs[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22296_ (.CLK(clknet_leaf_45_clk),
    .D(_01329_),
    .Q(\core.cpuregs[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22297_ (.CLK(clknet_leaf_71_clk),
    .D(_01330_),
    .Q(\core.cpuregs[31][19] ));
 sky130_fd_sc_hd__dfxtp_2 _22298_ (.CLK(clknet_leaf_53_clk),
    .D(_01331_),
    .Q(\core.cpuregs[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22299_ (.CLK(clknet_leaf_56_clk),
    .D(_01332_),
    .Q(\core.cpuregs[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22300_ (.CLK(clknet_leaf_61_clk),
    .D(_01333_),
    .Q(\core.cpuregs[31][22] ));
 sky130_fd_sc_hd__dfxtp_2 _22301_ (.CLK(clknet_leaf_53_clk),
    .D(_01334_),
    .Q(\core.cpuregs[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22302_ (.CLK(clknet_leaf_53_clk),
    .D(_01335_),
    .Q(\core.cpuregs[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22303_ (.CLK(clknet_leaf_58_clk),
    .D(_01336_),
    .Q(\core.cpuregs[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22304_ (.CLK(clknet_leaf_58_clk),
    .D(_01337_),
    .Q(\core.cpuregs[31][26] ));
 sky130_fd_sc_hd__dfxtp_2 _22305_ (.CLK(clknet_leaf_62_clk),
    .D(_01338_),
    .Q(\core.cpuregs[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22306_ (.CLK(clknet_leaf_62_clk),
    .D(_01339_),
    .Q(\core.cpuregs[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22307_ (.CLK(clknet_leaf_57_clk),
    .D(_01340_),
    .Q(\core.cpuregs[31][29] ));
 sky130_fd_sc_hd__dfxtp_2 _22308_ (.CLK(clknet_leaf_62_clk),
    .D(_01341_),
    .Q(\core.cpuregs[31][30] ));
 sky130_fd_sc_hd__dfxtp_2 _22309_ (.CLK(clknet_leaf_69_clk),
    .D(_01342_),
    .Q(\core.cpuregs[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22310_ (.CLK(clknet_leaf_25_clk),
    .D(_01343_),
    .Q(\core.mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22311_ (.CLK(clknet_leaf_37_clk),
    .D(_01344_),
    .Q(\core.mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22312_ (.CLK(clknet_leaf_3_clk),
    .D(_01345_),
    .Q(\core.mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22313_ (.CLK(clknet_leaf_79_clk),
    .D(_01346_),
    .Q(\core.mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22314_ (.CLK(clknet_leaf_5_clk),
    .D(_01347_),
    .Q(\core.mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22315_ (.CLK(clknet_leaf_4_clk),
    .D(_01348_),
    .Q(\core.mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22316_ (.CLK(clknet_leaf_4_clk),
    .D(_01349_),
    .Q(\core.mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _22317_ (.CLK(clknet_leaf_1_clk),
    .D(_01350_),
    .Q(\core.mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22318_ (.CLK(clknet_leaf_37_clk),
    .D(_01351_),
    .Q(\core.mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22319_ (.CLK(clknet_leaf_25_clk),
    .D(_01352_),
    .Q(\core.mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22320_ (.CLK(clknet_leaf_25_clk),
    .D(_01353_),
    .Q(\core.mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22321_ (.CLK(clknet_leaf_25_clk),
    .D(_01354_),
    .Q(\core.mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _22322_ (.CLK(clknet_leaf_25_clk),
    .D(_01355_),
    .Q(\core.mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _22323_ (.CLK(clknet_leaf_20_clk),
    .D(_01356_),
    .Q(\core.mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _22324_ (.CLK(clknet_leaf_21_clk),
    .D(_01357_),
    .Q(\core.mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _22325_ (.CLK(clknet_leaf_20_clk),
    .D(_01358_),
    .Q(\core.mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _22326_ (.CLK(clknet_leaf_25_clk),
    .D(_01359_),
    .Q(\core.mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _22327_ (.CLK(clknet_leaf_25_clk),
    .D(_01360_),
    .Q(\core.mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _22328_ (.CLK(clknet_leaf_2_clk),
    .D(_01361_),
    .Q(\core.mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _22329_ (.CLK(clknet_leaf_25_clk),
    .D(_01362_),
    .Q(\core.mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _22330_ (.CLK(clknet_leaf_20_clk),
    .D(_01363_),
    .Q(\core.mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _22331_ (.CLK(clknet_leaf_5_clk),
    .D(_01364_),
    .Q(\core.mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _22332_ (.CLK(clknet_leaf_17_clk),
    .D(_01365_),
    .Q(\core.mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _22333_ (.CLK(clknet_leaf_24_clk),
    .D(_01366_),
    .Q(\core.mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _22334_ (.CLK(clknet_leaf_20_clk),
    .D(_01367_),
    .Q(\core.mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _22335_ (.CLK(clknet_leaf_25_clk),
    .D(_01368_),
    .Q(\core.mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _22336_ (.CLK(clknet_leaf_24_clk),
    .D(_01369_),
    .Q(\core.mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _22337_ (.CLK(clknet_leaf_2_clk),
    .D(_01370_),
    .Q(\core.mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _22338_ (.CLK(clknet_leaf_23_clk),
    .D(_01371_),
    .Q(\core.mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _22339_ (.CLK(clknet_leaf_5_clk),
    .D(_01372_),
    .Q(\core.mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _22340_ (.CLK(clknet_leaf_2_clk),
    .D(_01373_),
    .Q(\core.mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _22341_ (.CLK(clknet_leaf_19_clk),
    .D(_01374_),
    .Q(\core.mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _22342_ (.CLK(clknet_leaf_37_clk),
    .D(_00025_),
    .Q(_00005_));
 sky130_fd_sc_hd__dfxtp_1 _22343_ (.CLK(clknet_leaf_37_clk),
    .D(_00026_),
    .Q(_00006_));
 sky130_fd_sc_hd__dfxtp_1 _22344_ (.CLK(clknet_leaf_37_clk),
    .D(_00027_),
    .Q(_00007_));
 sky130_fd_sc_hd__dfxtp_4 _22345_ (.CLK(clknet_leaf_79_clk),
    .D(_00028_),
    .Q(_00008_));
 sky130_fd_sc_hd__dfxtp_2 _22346_ (.CLK(clknet_leaf_37_clk),
    .D(_00029_),
    .Q(_00009_));
 sky130_fd_sc_hd__dfxtp_1 _22347_ (.CLK(clknet_leaf_45_clk),
    .D(_01375_),
    .Q(\core.cpuregs[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22348_ (.CLK(clknet_leaf_46_clk),
    .D(_01376_),
    .Q(\core.cpuregs[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22349_ (.CLK(clknet_leaf_85_clk),
    .D(_01377_),
    .Q(\core.cpuregs[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22350_ (.CLK(clknet_leaf_84_clk),
    .D(_01378_),
    .Q(\core.cpuregs[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22351_ (.CLK(clknet_leaf_84_clk),
    .D(_01379_),
    .Q(\core.cpuregs[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22352_ (.CLK(clknet_leaf_74_clk),
    .D(_01380_),
    .Q(\core.cpuregs[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22353_ (.CLK(clknet_leaf_75_clk),
    .D(_01381_),
    .Q(\core.cpuregs[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22354_ (.CLK(clknet_leaf_81_clk),
    .D(_01382_),
    .Q(\core.cpuregs[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22355_ (.CLK(clknet_leaf_69_clk),
    .D(_01383_),
    .Q(\core.cpuregs[29][8] ));
 sky130_fd_sc_hd__dfxtp_2 _22356_ (.CLK(clknet_leaf_67_clk),
    .D(_01384_),
    .Q(\core.cpuregs[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22357_ (.CLK(clknet_leaf_68_clk),
    .D(_01385_),
    .Q(\core.cpuregs[29][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22358_ (.CLK(clknet_leaf_46_clk),
    .D(_01386_),
    .Q(\core.cpuregs[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22359_ (.CLK(clknet_leaf_74_clk),
    .D(_01387_),
    .Q(\core.cpuregs[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22360_ (.CLK(clknet_leaf_46_clk),
    .D(_01388_),
    .Q(\core.cpuregs[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 _22361_ (.CLK(clknet_leaf_43_clk),
    .D(_01389_),
    .Q(\core.cpuregs[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 _22362_ (.CLK(clknet_leaf_72_clk),
    .D(_01390_),
    .Q(\core.cpuregs[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22363_ (.CLK(clknet_leaf_74_clk),
    .D(_01391_),
    .Q(\core.cpuregs[29][16] ));
 sky130_fd_sc_hd__dfxtp_2 _22364_ (.CLK(clknet_leaf_47_clk),
    .D(_01392_),
    .Q(\core.cpuregs[29][17] ));
 sky130_fd_sc_hd__dfxtp_2 _22365_ (.CLK(clknet_leaf_46_clk),
    .D(_01393_),
    .Q(\core.cpuregs[29][18] ));
 sky130_fd_sc_hd__dfxtp_2 _22366_ (.CLK(clknet_leaf_52_clk),
    .D(_01394_),
    .Q(\core.cpuregs[29][19] ));
 sky130_fd_sc_hd__dfxtp_2 _22367_ (.CLK(clknet_leaf_52_clk),
    .D(_01395_),
    .Q(\core.cpuregs[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22368_ (.CLK(clknet_leaf_55_clk),
    .D(_01396_),
    .Q(\core.cpuregs[29][21] ));
 sky130_fd_sc_hd__dfxtp_2 _22369_ (.CLK(clknet_leaf_70_clk),
    .D(_01397_),
    .Q(\core.cpuregs[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22370_ (.CLK(clknet_leaf_53_clk),
    .D(_01398_),
    .Q(\core.cpuregs[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22371_ (.CLK(clknet_leaf_55_clk),
    .D(_01399_),
    .Q(\core.cpuregs[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22372_ (.CLK(clknet_leaf_54_clk),
    .D(_01400_),
    .Q(\core.cpuregs[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22373_ (.CLK(clknet_leaf_58_clk),
    .D(_01401_),
    .Q(\core.cpuregs[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22374_ (.CLK(clknet_leaf_58_clk),
    .D(_01402_),
    .Q(\core.cpuregs[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22375_ (.CLK(clknet_leaf_63_clk),
    .D(_01403_),
    .Q(\core.cpuregs[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22376_ (.CLK(clknet_leaf_56_clk),
    .D(_01404_),
    .Q(\core.cpuregs[29][29] ));
 sky130_fd_sc_hd__dfxtp_2 _22377_ (.CLK(clknet_leaf_63_clk),
    .D(_01405_),
    .Q(\core.cpuregs[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22378_ (.CLK(clknet_leaf_70_clk),
    .D(_01406_),
    .Q(\core.cpuregs[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22379_ (.CLK(clknet_leaf_46_clk),
    .D(_01407_),
    .Q(\core.cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22380_ (.CLK(clknet_leaf_70_clk),
    .D(_01408_),
    .Q(\core.cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22381_ (.CLK(clknet_leaf_83_clk),
    .D(_01409_),
    .Q(\core.cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22382_ (.CLK(clknet_leaf_84_clk),
    .D(_01410_),
    .Q(\core.cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22383_ (.CLK(clknet_leaf_84_clk),
    .D(_01411_),
    .Q(\core.cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22384_ (.CLK(clknet_leaf_67_clk),
    .D(_01412_),
    .Q(\core.cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22385_ (.CLK(clknet_leaf_75_clk),
    .D(_01413_),
    .Q(\core.cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22386_ (.CLK(clknet_leaf_74_clk),
    .D(_01414_),
    .Q(\core.cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22387_ (.CLK(clknet_leaf_70_clk),
    .D(_01415_),
    .Q(\core.cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22388_ (.CLK(clknet_leaf_74_clk),
    .D(_01416_),
    .Q(\core.cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22389_ (.CLK(clknet_leaf_68_clk),
    .D(_01417_),
    .Q(\core.cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22390_ (.CLK(clknet_leaf_44_clk),
    .D(_01418_),
    .Q(\core.cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22391_ (.CLK(clknet_leaf_71_clk),
    .D(_01419_),
    .Q(\core.cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _22392_ (.CLK(clknet_leaf_45_clk),
    .D(_01420_),
    .Q(\core.cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _22393_ (.CLK(clknet_leaf_73_clk),
    .D(_01421_),
    .Q(\core.cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22394_ (.CLK(clknet_leaf_73_clk),
    .D(_01422_),
    .Q(\core.cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22395_ (.CLK(clknet_leaf_73_clk),
    .D(_01423_),
    .Q(\core.cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _22396_ (.CLK(clknet_leaf_43_clk),
    .D(_01424_),
    .Q(\core.cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22397_ (.CLK(clknet_leaf_46_clk),
    .D(_01425_),
    .Q(\core.cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _22398_ (.CLK(clknet_leaf_52_clk),
    .D(_01426_),
    .Q(\core.cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _22399_ (.CLK(clknet_leaf_52_clk),
    .D(_01427_),
    .Q(\core.cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22400_ (.CLK(clknet_leaf_56_clk),
    .D(_01428_),
    .Q(\core.cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22401_ (.CLK(clknet_leaf_57_clk),
    .D(_01429_),
    .Q(\core.cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22402_ (.CLK(clknet_leaf_55_clk),
    .D(_01430_),
    .Q(\core.cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22403_ (.CLK(clknet_leaf_55_clk),
    .D(_01431_),
    .Q(\core.cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22404_ (.CLK(clknet_leaf_56_clk),
    .D(_01432_),
    .Q(\core.cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22405_ (.CLK(clknet_leaf_62_clk),
    .D(_01433_),
    .Q(\core.cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22406_ (.CLK(clknet_leaf_62_clk),
    .D(_01434_),
    .Q(\core.cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22407_ (.CLK(clknet_leaf_62_clk),
    .D(_01435_),
    .Q(\core.cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22408_ (.CLK(clknet_leaf_58_clk),
    .D(_01436_),
    .Q(\core.cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _22409_ (.CLK(clknet_leaf_58_clk),
    .D(_01437_),
    .Q(\core.cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _22410_ (.CLK(clknet_leaf_70_clk),
    .D(_01438_),
    .Q(\core.cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22411_ (.CLK(clknet_leaf_68_clk),
    .D(_01439_),
    .Q(\core.cpuregs[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _22412_ (.CLK(clknet_leaf_71_clk),
    .D(_01440_),
    .Q(\core.cpuregs[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22413_ (.CLK(clknet_leaf_85_clk),
    .D(_01441_),
    .Q(\core.cpuregs[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _22414_ (.CLK(clknet_leaf_82_clk),
    .D(_01442_),
    .Q(\core.cpuregs[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22415_ (.CLK(clknet_leaf_83_clk),
    .D(_01443_),
    .Q(\core.cpuregs[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22416_ (.CLK(clknet_leaf_85_clk),
    .D(_01444_),
    .Q(\core.cpuregs[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _22417_ (.CLK(clknet_leaf_82_clk),
    .D(_01445_),
    .Q(\core.cpuregs[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22418_ (.CLK(clknet_leaf_82_clk),
    .D(_01446_),
    .Q(\core.cpuregs[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _22419_ (.CLK(clknet_leaf_70_clk),
    .D(_01447_),
    .Q(\core.cpuregs[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22420_ (.CLK(clknet_leaf_75_clk),
    .D(_01448_),
    .Q(\core.cpuregs[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22421_ (.CLK(clknet_leaf_72_clk),
    .D(_01449_),
    .Q(\core.cpuregs[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _22422_ (.CLK(clknet_leaf_45_clk),
    .D(_01450_),
    .Q(\core.cpuregs[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22423_ (.CLK(clknet_leaf_74_clk),
    .D(_01451_),
    .Q(\core.cpuregs[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22424_ (.CLK(clknet_leaf_44_clk),
    .D(_01452_),
    .Q(\core.cpuregs[24][13] ));
 sky130_fd_sc_hd__dfxtp_2 _22425_ (.CLK(clknet_leaf_73_clk),
    .D(_01453_),
    .Q(\core.cpuregs[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22426_ (.CLK(clknet_leaf_73_clk),
    .D(_01454_),
    .Q(\core.cpuregs[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22427_ (.CLK(clknet_leaf_76_clk),
    .D(_01455_),
    .Q(\core.cpuregs[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _22428_ (.CLK(clknet_leaf_43_clk),
    .D(_01456_),
    .Q(\core.cpuregs[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22429_ (.CLK(clknet_leaf_47_clk),
    .D(_01457_),
    .Q(\core.cpuregs[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _22430_ (.CLK(clknet_leaf_52_clk),
    .D(_01458_),
    .Q(\core.cpuregs[24][19] ));
 sky130_fd_sc_hd__dfxtp_2 _22431_ (.CLK(clknet_leaf_46_clk),
    .D(_01459_),
    .Q(\core.cpuregs[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22432_ (.CLK(clknet_leaf_53_clk),
    .D(_01460_),
    .Q(\core.cpuregs[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22433_ (.CLK(clknet_leaf_70_clk),
    .D(_01461_),
    .Q(\core.cpuregs[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22434_ (.CLK(clknet_leaf_57_clk),
    .D(_01462_),
    .Q(\core.cpuregs[24][23] ));
 sky130_fd_sc_hd__dfxtp_2 _22435_ (.CLK(clknet_leaf_52_clk),
    .D(_01463_),
    .Q(\core.cpuregs[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22436_ (.CLK(clknet_leaf_57_clk),
    .D(_01464_),
    .Q(\core.cpuregs[24][25] ));
 sky130_fd_sc_hd__dfxtp_2 _22437_ (.CLK(clknet_leaf_55_clk),
    .D(_01465_),
    .Q(\core.cpuregs[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22438_ (.CLK(clknet_leaf_62_clk),
    .D(_01466_),
    .Q(\core.cpuregs[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22439_ (.CLK(clknet_leaf_69_clk),
    .D(_01467_),
    .Q(\core.cpuregs[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22440_ (.CLK(clknet_leaf_69_clk),
    .D(_01468_),
    .Q(\core.cpuregs[24][29] ));
 sky130_fd_sc_hd__dfxtp_2 _22441_ (.CLK(clknet_leaf_62_clk),
    .D(_01469_),
    .Q(\core.cpuregs[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22442_ (.CLK(clknet_leaf_44_clk),
    .D(_01470_),
    .Q(\core.cpuregs[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22443_ (.CLK(clknet_leaf_39_clk),
    .D(_01471_),
    .Q(\core.cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _22444_ (.CLK(clknet_leaf_77_clk),
    .D(_01472_),
    .Q(\core.cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _22445_ (.CLK(clknet_leaf_82_clk),
    .D(_01473_),
    .Q(\core.cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _22446_ (.CLK(clknet_leaf_80_clk),
    .D(_01474_),
    .Q(\core.cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _22447_ (.CLK(clknet_leaf_83_clk),
    .D(_01475_),
    .Q(\core.cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _22448_ (.CLK(clknet_leaf_80_clk),
    .D(_01476_),
    .Q(\core.cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _22449_ (.CLK(clknet_leaf_80_clk),
    .D(_01477_),
    .Q(\core.cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _22450_ (.CLK(clknet_leaf_80_clk),
    .D(_01478_),
    .Q(\core.cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _22451_ (.CLK(clknet_leaf_76_clk),
    .D(_01479_),
    .Q(\core.cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _22452_ (.CLK(clknet_leaf_79_clk),
    .D(_01480_),
    .Q(\core.cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _22453_ (.CLK(clknet_leaf_78_clk),
    .D(_01481_),
    .Q(\core.cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _22454_ (.CLK(clknet_leaf_40_clk),
    .D(_01482_),
    .Q(\core.cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _22455_ (.CLK(clknet_leaf_78_clk),
    .D(_01483_),
    .Q(\core.cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _22456_ (.CLK(clknet_leaf_40_clk),
    .D(_01484_),
    .Q(\core.cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _22457_ (.CLK(clknet_leaf_38_clk),
    .D(_01485_),
    .Q(\core.cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _22458_ (.CLK(clknet_leaf_37_clk),
    .D(_01486_),
    .Q(\core.cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _22459_ (.CLK(clknet_leaf_37_clk),
    .D(_01487_),
    .Q(\core.cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _22460_ (.CLK(clknet_leaf_38_clk),
    .D(_01488_),
    .Q(\core.cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _22461_ (.CLK(clknet_leaf_41_clk),
    .D(_01489_),
    .Q(\core.cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _22462_ (.CLK(clknet_leaf_48_clk),
    .D(_01490_),
    .Q(\core.cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _22463_ (.CLK(clknet_leaf_40_clk),
    .D(_01491_),
    .Q(\core.cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _22464_ (.CLK(clknet_leaf_48_clk),
    .D(_01492_),
    .Q(\core.cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _22465_ (.CLK(clknet_leaf_48_clk),
    .D(_01493_),
    .Q(\core.cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _22466_ (.CLK(clknet_leaf_48_clk),
    .D(_01494_),
    .Q(\core.cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _22467_ (.CLK(clknet_leaf_41_clk),
    .D(_01495_),
    .Q(\core.cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _22468_ (.CLK(clknet_leaf_41_clk),
    .D(_01496_),
    .Q(\core.cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _22469_ (.CLK(clknet_leaf_48_clk),
    .D(_01497_),
    .Q(\core.cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _22470_ (.CLK(clknet_leaf_48_clk),
    .D(_01498_),
    .Q(\core.cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _22471_ (.CLK(clknet_leaf_78_clk),
    .D(_01499_),
    .Q(\core.cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _22472_ (.CLK(clknet_leaf_35_clk),
    .D(_01500_),
    .Q(\core.cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _22473_ (.CLK(clknet_leaf_48_clk),
    .D(_01501_),
    .Q(\core.cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _22474_ (.CLK(clknet_leaf_41_clk),
    .D(_01502_),
    .Q(\core.cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _22475_ (.CLK(clknet_leaf_6_clk),
    .D(_01503_),
    .Q(\core.instr_lhu ));
 sky130_fd_sc_hd__dfxtp_1 _22476_ (.CLK(clknet_leaf_17_clk),
    .D(_01504_),
    .Q(\core.instr_lbu ));
 sky130_fd_sc_hd__dfxtp_1 _22477_ (.CLK(clknet_leaf_17_clk),
    .D(_01505_),
    .Q(\core.instr_lw ));
 sky130_fd_sc_hd__dfxtp_1 _22478_ (.CLK(clknet_leaf_6_clk),
    .D(_01506_),
    .Q(\core.instr_lh ));
 sky130_fd_sc_hd__dfxtp_1 _22479_ (.CLK(clknet_leaf_6_clk),
    .D(_01507_),
    .Q(\core.instr_bgeu ));
 sky130_fd_sc_hd__dfxtp_1 _22480_ (.CLK(clknet_leaf_6_clk),
    .D(_01508_),
    .Q(\core.instr_blt ));
 sky130_fd_sc_hd__dfxtp_2 _22481_ (.CLK(clknet_leaf_2_clk),
    .D(_00034_),
    .Q(\core.reg_sh[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22482_ (.CLK(clknet_leaf_24_clk),
    .D(_00035_),
    .Q(\core.reg_sh[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22483_ (.CLK(clknet_leaf_2_clk),
    .D(_00036_),
    .Q(\core.reg_sh[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22484_ (.CLK(clknet_leaf_19_clk),
    .D(_01509_),
    .Q(\core.instr_rdinstrh ));
 sky130_fd_sc_hd__dfxtp_1 _22485_ (.CLK(clknet_leaf_37_clk),
    .D(_00020_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_2 _22486_ (.CLK(clknet_leaf_78_clk),
    .D(_00021_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_1 _22487_ (.CLK(clknet_leaf_79_clk),
    .D(_00022_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_2 _22488_ (.CLK(clknet_leaf_78_clk),
    .D(_00023_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_1 _22489_ (.CLK(clknet_leaf_37_clk),
    .D(_00024_),
    .Q(_00004_));
 sky130_fd_sc_hd__dfxtp_1 _22490_ (.CLK(clknet_leaf_19_clk),
    .D(_01510_),
    .Q(\core.instr_rdinstr ));
 sky130_fd_sc_hd__dfxtp_1 _22491_ (.CLK(clknet_leaf_6_clk),
    .D(_01511_),
    .Q(\core.instr_rdcycle ));
 sky130_fd_sc_hd__dfxtp_1 _22492_ (.CLK(clknet_leaf_6_clk),
    .D(_01512_),
    .Q(\core.instr_srai ));
 sky130_fd_sc_hd__dfxtp_1 _22493_ (.CLK(clknet_leaf_6_clk),
    .D(_01513_),
    .Q(\core.instr_and ));
 sky130_fd_sc_hd__dfxtp_1 _22494_ (.CLK(clknet_leaf_17_clk),
    .D(_01514_),
    .Q(\core.instr_or ));
 sky130_fd_sc_hd__dfxtp_1 _22495_ (.CLK(clknet_leaf_6_clk),
    .D(_01515_),
    .Q(\core.instr_srl ));
 sky130_fd_sc_hd__dfxtp_1 _22496_ (.CLK(clknet_leaf_17_clk),
    .D(_01516_),
    .Q(\core.instr_sltu ));
 sky130_fd_sc_hd__dfxtp_1 _22497_ (.CLK(clknet_leaf_17_clk),
    .D(_01517_),
    .Q(\core.instr_slt ));
 sky130_fd_sc_hd__dfxtp_1 _22498_ (.CLK(clknet_leaf_5_clk),
    .D(_01518_),
    .Q(\core.instr_sub ));
 sky130_fd_sc_hd__dfxtp_1 _22499_ (.CLK(clknet_leaf_17_clk),
    .D(_01519_),
    .Q(\core.instr_slli ));
 sky130_fd_sc_hd__dfxtp_1 _22500_ (.CLK(clknet_leaf_18_clk),
    .D(_01520_),
    .Q(\core.instr_sw ));
 sky130_fd_sc_hd__dfxtp_1 _22501_ (.CLK(clknet_leaf_17_clk),
    .D(_01521_),
    .Q(\core.instr_andi ));
 sky130_fd_sc_hd__dfxtp_1 _22502_ (.CLK(clknet_leaf_6_clk),
    .D(_01522_),
    .Q(\core.instr_xori ));
 sky130_fd_sc_hd__dfxtp_1 _22503_ (.CLK(clknet_leaf_6_clk),
    .D(_01523_),
    .Q(\core.instr_addi ));
 sky130_fd_sc_hd__dfxtp_1 _22504_ (.CLK(clknet_leaf_19_clk),
    .D(_01524_),
    .Q(\core.instr_sb ));
 sky130_fd_sc_hd__dfxtp_1 _22505_ (.CLK(clknet_leaf_24_clk),
    .D(_01525_),
    .Q(\core.mem_do_rdata ));
 sky130_fd_sc_hd__dfxtp_1 _22506_ (.CLK(clknet_leaf_24_clk),
    .D(_01526_),
    .Q(\core.mem_do_rinst ));
 sky130_fd_sc_hd__dfxtp_1 _22507_ (.CLK(clknet_leaf_22_clk),
    .D(_01527_),
    .Q(\core.mem_do_prefetch ));
 sky130_fd_sc_hd__dfxtp_1 _22508_ (.CLK(clknet_leaf_87_clk),
    .D(_01528_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_2 _22509_ (.CLK(clknet_leaf_27_clk),
    .D(_01529_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _22510_ (.CLK(clknet_leaf_8_clk),
    .D(_01530_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _22511_ (.CLK(clknet_leaf_88_clk),
    .D(_01531_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_2 _22512_ (.CLK(clknet_leaf_90_clk),
    .D(_01532_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _22513_ (.CLK(clknet_leaf_29_clk),
    .D(_01533_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _22514_ (.CLK(clknet_leaf_89_clk),
    .D(_01534_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_2 _22515_ (.CLK(clknet_leaf_91_clk),
    .D(_01535_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_2 _22516_ (.CLK(clknet_3_7__leaf_clk),
    .D(_01536_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _22517_ (.CLK(clknet_leaf_7_clk),
    .D(_01537_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _22518_ (.CLK(clknet_leaf_8_clk),
    .D(_01538_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _22519_ (.CLK(clknet_leaf_27_clk),
    .D(_01539_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _22520_ (.CLK(clknet_leaf_28_clk),
    .D(_01540_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _22521_ (.CLK(clknet_leaf_91_clk),
    .D(_01541_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _22522_ (.CLK(clknet_leaf_7_clk),
    .D(_01542_),
    .Q(net41));
 sky130_fd_sc_hd__conb_1 picorv32_wrapper_107 (.LO(net107));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(mem_rdata[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(mem_rdata[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(mem_rdata[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(mem_rdata[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(mem_rdata[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(mem_rdata[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(mem_rdata[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(mem_rdata[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(mem_rdata[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(mem_rdata[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(mem_rdata[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(mem_rdata[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(mem_rdata[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(mem_rdata[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(mem_rdata[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(mem_rdata[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(mem_rdata[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(mem_rdata[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(mem_rdata[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(mem_rdata[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(mem_rdata[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(mem_rdata[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(mem_rdata[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(mem_rdata[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(mem_rdata[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(mem_rdata[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(mem_rdata[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(mem_rdata[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(mem_rdata[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(mem_rdata[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(mem_rdata[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(mem_rdata[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(mem_ready),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(resetn),
    .X(net34));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_4 output41 (.A(net41),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_4 output45 (.A(net45),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_4 output60 (.A(net60),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(mem_instr));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net87),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(trap));
 sky130_fd_sc_hd__clkbuf_2 max_cap104 (.A(_07009_),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap105 (.A(_07614_),
    .X(net105));
 sky130_fd_sc_hd__conb_1 picorv32_wrapper_106 (.LO(net106));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\core.mem_wordsize[0] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net100),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\core.instr_rdcycle ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\core.reg_next_pc[3] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\core.count_cycle[34] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\core.reg_next_pc[22] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net102),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net65),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\core.reg_next_pc[23] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\core.cpuregs[30][29] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net99),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\core.instr_slli ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\core.cpuregs[17][21] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\core.cpuregs[18][24] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\core.reg_next_pc[6] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\core.cpuregs[10][28] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\core.cpuregs[28][20] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\core.cpuregs[3][28] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\core.cpuregs[7][23] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\core.cpuregs[17][19] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\core.cpuregs[1][30] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\core.cpuregs[27][20] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\core.cpuregs[12][28] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\core.cpuregs[14][25] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\core.cpuregs[13][24] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\core.reg_next_pc[20] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\core.cpuregs[6][31] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\core.reg_next_pc[13] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_00129_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\core.cpuregs[12][26] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\core.cpuregs[29][21] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\core.cpuregs[14][31] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\core.cpuregs[10][31] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\core.cpuregs[12][19] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\core.cpuregs[14][26] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\core.cpuregs[8][26] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\core.cpuregs[12][24] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\core.cpuregs[1][21] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\core.cpuregs[8][23] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\core.cpuregs[31][19] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\core.cpuregs[10][24] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\core.cpuregs[8][24] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\core.cpuregs[9][30] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\core.cpuregs[6][30] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\core.cpuregs[22][31] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\core.cpuregs[28][29] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\core.cpuregs[9][24] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\core.cpuregs[8][30] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\core.cpuregs[10][23] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\core.cpuregs[4][31] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\core.cpuregs[27][22] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\core.cpuregs[15][19] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\core.cpuregs[13][21] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\core.cpuregs[2][19] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\core.cpuregs[2][23] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\core.cpuregs[5][23] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\core.cpuregs[18][21] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\core.cpuregs[8][21] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\core.cpuregs[4][24] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\core.cpuregs[13][22] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\core.cpuregs[9][21] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\core.cpuregs[24][31] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\core.cpuregs[12][29] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\core.cpuregs[9][23] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\core.cpuregs[4][23] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\core.cpuregs[10][27] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\core.cpuregs[10][22] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\core.cpuregs[28][31] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\core.is_compare ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\core.cpuregs[24][21] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\core.cpuregs[5][31] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\core.cpuregs[2][25] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\core.cpuregs[3][21] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\core.cpuregs[24][20] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\core.cpuregs[9][28] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\core.cpuregs[11][27] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\core.cpuregs[18][27] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\core.cpuregs[27][23] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\core.cpuregs[4][22] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\core.cpuregs[7][26] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\core.reg_next_pc[24] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\core.cpuregs[2][31] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\core.cpuregs[21][30] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\core.cpuregs[9][29] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\core.reg_sh[1] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\core.cpuregs[2][21] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\core.cpuregs[15][21] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\core.cpuregs[20][26] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\core.cpuregs[27][19] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\core.cpuregs[6][25] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\core.cpuregs[28][19] ),
    .X(net198));
 assign mem_addr[0] = net106;
 assign mem_addr[1] = net107;
endmodule
