module picorv32_wrapper (clk,
    mem_instr,
    mem_ready,
    mem_valid,
    resetn,
    trap,
    mem_addr,
    mem_rdata,
    mem_wdata,
    mem_wstrb);
 input clk;
 output mem_instr;
 input mem_ready;
 output mem_valid;
 input resetn;
 output trap;
 output [31:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire \core.alu_out[0] ;
 wire \core.alu_out[10] ;
 wire \core.alu_out[11] ;
 wire \core.alu_out[12] ;
 wire \core.alu_out[13] ;
 wire \core.alu_out[14] ;
 wire \core.alu_out[15] ;
 wire \core.alu_out[16] ;
 wire \core.alu_out[17] ;
 wire \core.alu_out[18] ;
 wire \core.alu_out[19] ;
 wire \core.alu_out[1] ;
 wire \core.alu_out[20] ;
 wire \core.alu_out[21] ;
 wire \core.alu_out[22] ;
 wire \core.alu_out[23] ;
 wire \core.alu_out[24] ;
 wire \core.alu_out[25] ;
 wire \core.alu_out[26] ;
 wire \core.alu_out[27] ;
 wire \core.alu_out[28] ;
 wire \core.alu_out[29] ;
 wire \core.alu_out[2] ;
 wire \core.alu_out[30] ;
 wire \core.alu_out[31] ;
 wire \core.alu_out[3] ;
 wire \core.alu_out[4] ;
 wire \core.alu_out[5] ;
 wire \core.alu_out[6] ;
 wire \core.alu_out[7] ;
 wire \core.alu_out[8] ;
 wire \core.alu_out[9] ;
 wire \core.alu_out_q[0] ;
 wire \core.alu_out_q[10] ;
 wire \core.alu_out_q[11] ;
 wire \core.alu_out_q[12] ;
 wire \core.alu_out_q[13] ;
 wire \core.alu_out_q[14] ;
 wire \core.alu_out_q[15] ;
 wire \core.alu_out_q[16] ;
 wire \core.alu_out_q[17] ;
 wire \core.alu_out_q[18] ;
 wire \core.alu_out_q[19] ;
 wire \core.alu_out_q[1] ;
 wire \core.alu_out_q[20] ;
 wire \core.alu_out_q[21] ;
 wire \core.alu_out_q[22] ;
 wire \core.alu_out_q[23] ;
 wire \core.alu_out_q[24] ;
 wire \core.alu_out_q[25] ;
 wire \core.alu_out_q[26] ;
 wire \core.alu_out_q[27] ;
 wire \core.alu_out_q[28] ;
 wire \core.alu_out_q[29] ;
 wire \core.alu_out_q[2] ;
 wire \core.alu_out_q[30] ;
 wire \core.alu_out_q[31] ;
 wire \core.alu_out_q[3] ;
 wire \core.alu_out_q[4] ;
 wire \core.alu_out_q[5] ;
 wire \core.alu_out_q[6] ;
 wire \core.alu_out_q[7] ;
 wire \core.alu_out_q[8] ;
 wire \core.alu_out_q[9] ;
 wire \core.count_cycle[0] ;
 wire \core.count_cycle[10] ;
 wire \core.count_cycle[11] ;
 wire \core.count_cycle[12] ;
 wire \core.count_cycle[13] ;
 wire \core.count_cycle[14] ;
 wire \core.count_cycle[15] ;
 wire \core.count_cycle[16] ;
 wire \core.count_cycle[17] ;
 wire \core.count_cycle[18] ;
 wire \core.count_cycle[19] ;
 wire \core.count_cycle[1] ;
 wire \core.count_cycle[20] ;
 wire \core.count_cycle[21] ;
 wire \core.count_cycle[22] ;
 wire \core.count_cycle[23] ;
 wire \core.count_cycle[24] ;
 wire \core.count_cycle[25] ;
 wire \core.count_cycle[26] ;
 wire \core.count_cycle[27] ;
 wire \core.count_cycle[28] ;
 wire \core.count_cycle[29] ;
 wire \core.count_cycle[2] ;
 wire \core.count_cycle[30] ;
 wire \core.count_cycle[31] ;
 wire \core.count_cycle[32] ;
 wire \core.count_cycle[33] ;
 wire \core.count_cycle[34] ;
 wire \core.count_cycle[35] ;
 wire \core.count_cycle[36] ;
 wire \core.count_cycle[37] ;
 wire \core.count_cycle[38] ;
 wire \core.count_cycle[39] ;
 wire \core.count_cycle[3] ;
 wire \core.count_cycle[40] ;
 wire \core.count_cycle[41] ;
 wire \core.count_cycle[42] ;
 wire \core.count_cycle[43] ;
 wire \core.count_cycle[44] ;
 wire \core.count_cycle[45] ;
 wire \core.count_cycle[46] ;
 wire \core.count_cycle[47] ;
 wire \core.count_cycle[48] ;
 wire \core.count_cycle[49] ;
 wire \core.count_cycle[4] ;
 wire \core.count_cycle[50] ;
 wire \core.count_cycle[51] ;
 wire \core.count_cycle[52] ;
 wire \core.count_cycle[53] ;
 wire \core.count_cycle[54] ;
 wire \core.count_cycle[55] ;
 wire \core.count_cycle[56] ;
 wire \core.count_cycle[57] ;
 wire \core.count_cycle[58] ;
 wire \core.count_cycle[59] ;
 wire \core.count_cycle[5] ;
 wire \core.count_cycle[60] ;
 wire \core.count_cycle[61] ;
 wire \core.count_cycle[62] ;
 wire \core.count_cycle[63] ;
 wire \core.count_cycle[6] ;
 wire \core.count_cycle[7] ;
 wire \core.count_cycle[8] ;
 wire \core.count_cycle[9] ;
 wire \core.count_instr[0] ;
 wire \core.count_instr[10] ;
 wire \core.count_instr[11] ;
 wire \core.count_instr[12] ;
 wire \core.count_instr[13] ;
 wire \core.count_instr[14] ;
 wire \core.count_instr[15] ;
 wire \core.count_instr[16] ;
 wire \core.count_instr[17] ;
 wire \core.count_instr[18] ;
 wire \core.count_instr[19] ;
 wire \core.count_instr[1] ;
 wire \core.count_instr[20] ;
 wire \core.count_instr[21] ;
 wire \core.count_instr[22] ;
 wire \core.count_instr[23] ;
 wire \core.count_instr[24] ;
 wire \core.count_instr[25] ;
 wire \core.count_instr[26] ;
 wire \core.count_instr[27] ;
 wire \core.count_instr[28] ;
 wire \core.count_instr[29] ;
 wire \core.count_instr[2] ;
 wire \core.count_instr[30] ;
 wire \core.count_instr[31] ;
 wire \core.count_instr[32] ;
 wire \core.count_instr[33] ;
 wire \core.count_instr[34] ;
 wire \core.count_instr[35] ;
 wire \core.count_instr[36] ;
 wire \core.count_instr[37] ;
 wire \core.count_instr[38] ;
 wire \core.count_instr[39] ;
 wire \core.count_instr[3] ;
 wire \core.count_instr[40] ;
 wire \core.count_instr[41] ;
 wire \core.count_instr[42] ;
 wire \core.count_instr[43] ;
 wire \core.count_instr[44] ;
 wire \core.count_instr[45] ;
 wire \core.count_instr[46] ;
 wire \core.count_instr[47] ;
 wire \core.count_instr[48] ;
 wire \core.count_instr[49] ;
 wire \core.count_instr[4] ;
 wire \core.count_instr[50] ;
 wire \core.count_instr[51] ;
 wire \core.count_instr[52] ;
 wire \core.count_instr[53] ;
 wire \core.count_instr[54] ;
 wire \core.count_instr[55] ;
 wire \core.count_instr[56] ;
 wire \core.count_instr[57] ;
 wire \core.count_instr[58] ;
 wire \core.count_instr[59] ;
 wire \core.count_instr[5] ;
 wire \core.count_instr[60] ;
 wire \core.count_instr[61] ;
 wire \core.count_instr[62] ;
 wire \core.count_instr[63] ;
 wire \core.count_instr[6] ;
 wire \core.count_instr[7] ;
 wire \core.count_instr[8] ;
 wire \core.count_instr[9] ;
 wire \core.cpu_state[0] ;
 wire \core.cpu_state[1] ;
 wire \core.cpu_state[2] ;
 wire \core.cpu_state[3] ;
 wire \core.cpu_state[4] ;
 wire \core.cpu_state[5] ;
 wire \core.cpu_state[6] ;
 wire \core.cpuregs[0][0] ;
 wire \core.cpuregs[0][10] ;
 wire \core.cpuregs[0][11] ;
 wire \core.cpuregs[0][12] ;
 wire \core.cpuregs[0][13] ;
 wire \core.cpuregs[0][14] ;
 wire \core.cpuregs[0][15] ;
 wire \core.cpuregs[0][16] ;
 wire \core.cpuregs[0][17] ;
 wire \core.cpuregs[0][18] ;
 wire \core.cpuregs[0][19] ;
 wire \core.cpuregs[0][1] ;
 wire \core.cpuregs[0][20] ;
 wire \core.cpuregs[0][21] ;
 wire \core.cpuregs[0][22] ;
 wire \core.cpuregs[0][23] ;
 wire \core.cpuregs[0][24] ;
 wire \core.cpuregs[0][25] ;
 wire \core.cpuregs[0][26] ;
 wire \core.cpuregs[0][27] ;
 wire \core.cpuregs[0][28] ;
 wire \core.cpuregs[0][29] ;
 wire \core.cpuregs[0][2] ;
 wire \core.cpuregs[0][30] ;
 wire \core.cpuregs[0][31] ;
 wire \core.cpuregs[0][3] ;
 wire \core.cpuregs[0][4] ;
 wire \core.cpuregs[0][5] ;
 wire \core.cpuregs[0][6] ;
 wire \core.cpuregs[0][7] ;
 wire \core.cpuregs[0][8] ;
 wire \core.cpuregs[0][9] ;
 wire \core.cpuregs[10][0] ;
 wire \core.cpuregs[10][10] ;
 wire \core.cpuregs[10][11] ;
 wire \core.cpuregs[10][12] ;
 wire \core.cpuregs[10][13] ;
 wire \core.cpuregs[10][14] ;
 wire \core.cpuregs[10][15] ;
 wire \core.cpuregs[10][16] ;
 wire \core.cpuregs[10][17] ;
 wire \core.cpuregs[10][18] ;
 wire \core.cpuregs[10][19] ;
 wire \core.cpuregs[10][1] ;
 wire \core.cpuregs[10][20] ;
 wire \core.cpuregs[10][21] ;
 wire \core.cpuregs[10][22] ;
 wire \core.cpuregs[10][23] ;
 wire \core.cpuregs[10][24] ;
 wire \core.cpuregs[10][25] ;
 wire \core.cpuregs[10][26] ;
 wire \core.cpuregs[10][27] ;
 wire \core.cpuregs[10][28] ;
 wire \core.cpuregs[10][29] ;
 wire \core.cpuregs[10][2] ;
 wire \core.cpuregs[10][30] ;
 wire \core.cpuregs[10][31] ;
 wire \core.cpuregs[10][3] ;
 wire \core.cpuregs[10][4] ;
 wire \core.cpuregs[10][5] ;
 wire \core.cpuregs[10][6] ;
 wire \core.cpuregs[10][7] ;
 wire \core.cpuregs[10][8] ;
 wire \core.cpuregs[10][9] ;
 wire \core.cpuregs[11][0] ;
 wire \core.cpuregs[11][10] ;
 wire \core.cpuregs[11][11] ;
 wire \core.cpuregs[11][12] ;
 wire \core.cpuregs[11][13] ;
 wire \core.cpuregs[11][14] ;
 wire \core.cpuregs[11][15] ;
 wire \core.cpuregs[11][16] ;
 wire \core.cpuregs[11][17] ;
 wire \core.cpuregs[11][18] ;
 wire \core.cpuregs[11][19] ;
 wire \core.cpuregs[11][1] ;
 wire \core.cpuregs[11][20] ;
 wire \core.cpuregs[11][21] ;
 wire \core.cpuregs[11][22] ;
 wire \core.cpuregs[11][23] ;
 wire \core.cpuregs[11][24] ;
 wire \core.cpuregs[11][25] ;
 wire \core.cpuregs[11][26] ;
 wire \core.cpuregs[11][27] ;
 wire \core.cpuregs[11][28] ;
 wire \core.cpuregs[11][29] ;
 wire \core.cpuregs[11][2] ;
 wire \core.cpuregs[11][30] ;
 wire \core.cpuregs[11][31] ;
 wire \core.cpuregs[11][3] ;
 wire \core.cpuregs[11][4] ;
 wire \core.cpuregs[11][5] ;
 wire \core.cpuregs[11][6] ;
 wire \core.cpuregs[11][7] ;
 wire \core.cpuregs[11][8] ;
 wire \core.cpuregs[11][9] ;
 wire \core.cpuregs[12][0] ;
 wire \core.cpuregs[12][10] ;
 wire \core.cpuregs[12][11] ;
 wire \core.cpuregs[12][12] ;
 wire \core.cpuregs[12][13] ;
 wire \core.cpuregs[12][14] ;
 wire \core.cpuregs[12][15] ;
 wire \core.cpuregs[12][16] ;
 wire \core.cpuregs[12][17] ;
 wire \core.cpuregs[12][18] ;
 wire \core.cpuregs[12][19] ;
 wire \core.cpuregs[12][1] ;
 wire \core.cpuregs[12][20] ;
 wire \core.cpuregs[12][21] ;
 wire \core.cpuregs[12][22] ;
 wire \core.cpuregs[12][23] ;
 wire \core.cpuregs[12][24] ;
 wire \core.cpuregs[12][25] ;
 wire \core.cpuregs[12][26] ;
 wire \core.cpuregs[12][27] ;
 wire \core.cpuregs[12][28] ;
 wire \core.cpuregs[12][29] ;
 wire \core.cpuregs[12][2] ;
 wire \core.cpuregs[12][30] ;
 wire \core.cpuregs[12][31] ;
 wire \core.cpuregs[12][3] ;
 wire \core.cpuregs[12][4] ;
 wire \core.cpuregs[12][5] ;
 wire \core.cpuregs[12][6] ;
 wire \core.cpuregs[12][7] ;
 wire \core.cpuregs[12][8] ;
 wire \core.cpuregs[12][9] ;
 wire \core.cpuregs[13][0] ;
 wire \core.cpuregs[13][10] ;
 wire \core.cpuregs[13][11] ;
 wire \core.cpuregs[13][12] ;
 wire \core.cpuregs[13][13] ;
 wire \core.cpuregs[13][14] ;
 wire \core.cpuregs[13][15] ;
 wire \core.cpuregs[13][16] ;
 wire \core.cpuregs[13][17] ;
 wire \core.cpuregs[13][18] ;
 wire \core.cpuregs[13][19] ;
 wire \core.cpuregs[13][1] ;
 wire \core.cpuregs[13][20] ;
 wire \core.cpuregs[13][21] ;
 wire \core.cpuregs[13][22] ;
 wire \core.cpuregs[13][23] ;
 wire \core.cpuregs[13][24] ;
 wire \core.cpuregs[13][25] ;
 wire \core.cpuregs[13][26] ;
 wire \core.cpuregs[13][27] ;
 wire \core.cpuregs[13][28] ;
 wire \core.cpuregs[13][29] ;
 wire \core.cpuregs[13][2] ;
 wire \core.cpuregs[13][30] ;
 wire \core.cpuregs[13][31] ;
 wire \core.cpuregs[13][3] ;
 wire \core.cpuregs[13][4] ;
 wire \core.cpuregs[13][5] ;
 wire \core.cpuregs[13][6] ;
 wire \core.cpuregs[13][7] ;
 wire \core.cpuregs[13][8] ;
 wire \core.cpuregs[13][9] ;
 wire \core.cpuregs[14][0] ;
 wire \core.cpuregs[14][10] ;
 wire \core.cpuregs[14][11] ;
 wire \core.cpuregs[14][12] ;
 wire \core.cpuregs[14][13] ;
 wire \core.cpuregs[14][14] ;
 wire \core.cpuregs[14][15] ;
 wire \core.cpuregs[14][16] ;
 wire \core.cpuregs[14][17] ;
 wire \core.cpuregs[14][18] ;
 wire \core.cpuregs[14][19] ;
 wire \core.cpuregs[14][1] ;
 wire \core.cpuregs[14][20] ;
 wire \core.cpuregs[14][21] ;
 wire \core.cpuregs[14][22] ;
 wire \core.cpuregs[14][23] ;
 wire \core.cpuregs[14][24] ;
 wire \core.cpuregs[14][25] ;
 wire \core.cpuregs[14][26] ;
 wire \core.cpuregs[14][27] ;
 wire \core.cpuregs[14][28] ;
 wire \core.cpuregs[14][29] ;
 wire \core.cpuregs[14][2] ;
 wire \core.cpuregs[14][30] ;
 wire \core.cpuregs[14][31] ;
 wire \core.cpuregs[14][3] ;
 wire \core.cpuregs[14][4] ;
 wire \core.cpuregs[14][5] ;
 wire \core.cpuregs[14][6] ;
 wire \core.cpuregs[14][7] ;
 wire \core.cpuregs[14][8] ;
 wire \core.cpuregs[14][9] ;
 wire \core.cpuregs[15][0] ;
 wire \core.cpuregs[15][10] ;
 wire \core.cpuregs[15][11] ;
 wire \core.cpuregs[15][12] ;
 wire \core.cpuregs[15][13] ;
 wire \core.cpuregs[15][14] ;
 wire \core.cpuregs[15][15] ;
 wire \core.cpuregs[15][16] ;
 wire \core.cpuregs[15][17] ;
 wire \core.cpuregs[15][18] ;
 wire \core.cpuregs[15][19] ;
 wire \core.cpuregs[15][1] ;
 wire \core.cpuregs[15][20] ;
 wire \core.cpuregs[15][21] ;
 wire \core.cpuregs[15][22] ;
 wire \core.cpuregs[15][23] ;
 wire \core.cpuregs[15][24] ;
 wire \core.cpuregs[15][25] ;
 wire \core.cpuregs[15][26] ;
 wire \core.cpuregs[15][27] ;
 wire \core.cpuregs[15][28] ;
 wire \core.cpuregs[15][29] ;
 wire \core.cpuregs[15][2] ;
 wire \core.cpuregs[15][30] ;
 wire \core.cpuregs[15][31] ;
 wire \core.cpuregs[15][3] ;
 wire \core.cpuregs[15][4] ;
 wire \core.cpuregs[15][5] ;
 wire \core.cpuregs[15][6] ;
 wire \core.cpuregs[15][7] ;
 wire \core.cpuregs[15][8] ;
 wire \core.cpuregs[15][9] ;
 wire \core.cpuregs[16][0] ;
 wire \core.cpuregs[16][10] ;
 wire \core.cpuregs[16][11] ;
 wire \core.cpuregs[16][12] ;
 wire \core.cpuregs[16][13] ;
 wire \core.cpuregs[16][14] ;
 wire \core.cpuregs[16][15] ;
 wire \core.cpuregs[16][16] ;
 wire \core.cpuregs[16][17] ;
 wire \core.cpuregs[16][18] ;
 wire \core.cpuregs[16][19] ;
 wire \core.cpuregs[16][1] ;
 wire \core.cpuregs[16][20] ;
 wire \core.cpuregs[16][21] ;
 wire \core.cpuregs[16][22] ;
 wire \core.cpuregs[16][23] ;
 wire \core.cpuregs[16][24] ;
 wire \core.cpuregs[16][25] ;
 wire \core.cpuregs[16][26] ;
 wire \core.cpuregs[16][27] ;
 wire \core.cpuregs[16][28] ;
 wire \core.cpuregs[16][29] ;
 wire \core.cpuregs[16][2] ;
 wire \core.cpuregs[16][30] ;
 wire \core.cpuregs[16][31] ;
 wire \core.cpuregs[16][3] ;
 wire \core.cpuregs[16][4] ;
 wire \core.cpuregs[16][5] ;
 wire \core.cpuregs[16][6] ;
 wire \core.cpuregs[16][7] ;
 wire \core.cpuregs[16][8] ;
 wire \core.cpuregs[16][9] ;
 wire \core.cpuregs[17][0] ;
 wire \core.cpuregs[17][10] ;
 wire \core.cpuregs[17][11] ;
 wire \core.cpuregs[17][12] ;
 wire \core.cpuregs[17][13] ;
 wire \core.cpuregs[17][14] ;
 wire \core.cpuregs[17][15] ;
 wire \core.cpuregs[17][16] ;
 wire \core.cpuregs[17][17] ;
 wire \core.cpuregs[17][18] ;
 wire \core.cpuregs[17][19] ;
 wire \core.cpuregs[17][1] ;
 wire \core.cpuregs[17][20] ;
 wire \core.cpuregs[17][21] ;
 wire \core.cpuregs[17][22] ;
 wire \core.cpuregs[17][23] ;
 wire \core.cpuregs[17][24] ;
 wire \core.cpuregs[17][25] ;
 wire \core.cpuregs[17][26] ;
 wire \core.cpuregs[17][27] ;
 wire \core.cpuregs[17][28] ;
 wire \core.cpuregs[17][29] ;
 wire \core.cpuregs[17][2] ;
 wire \core.cpuregs[17][30] ;
 wire \core.cpuregs[17][31] ;
 wire \core.cpuregs[17][3] ;
 wire \core.cpuregs[17][4] ;
 wire \core.cpuregs[17][5] ;
 wire \core.cpuregs[17][6] ;
 wire \core.cpuregs[17][7] ;
 wire \core.cpuregs[17][8] ;
 wire \core.cpuregs[17][9] ;
 wire \core.cpuregs[18][0] ;
 wire \core.cpuregs[18][10] ;
 wire \core.cpuregs[18][11] ;
 wire \core.cpuregs[18][12] ;
 wire \core.cpuregs[18][13] ;
 wire \core.cpuregs[18][14] ;
 wire \core.cpuregs[18][15] ;
 wire \core.cpuregs[18][16] ;
 wire \core.cpuregs[18][17] ;
 wire \core.cpuregs[18][18] ;
 wire \core.cpuregs[18][19] ;
 wire \core.cpuregs[18][1] ;
 wire \core.cpuregs[18][20] ;
 wire \core.cpuregs[18][21] ;
 wire \core.cpuregs[18][22] ;
 wire \core.cpuregs[18][23] ;
 wire \core.cpuregs[18][24] ;
 wire \core.cpuregs[18][25] ;
 wire \core.cpuregs[18][26] ;
 wire \core.cpuregs[18][27] ;
 wire \core.cpuregs[18][28] ;
 wire \core.cpuregs[18][29] ;
 wire \core.cpuregs[18][2] ;
 wire \core.cpuregs[18][30] ;
 wire \core.cpuregs[18][31] ;
 wire \core.cpuregs[18][3] ;
 wire \core.cpuregs[18][4] ;
 wire \core.cpuregs[18][5] ;
 wire \core.cpuregs[18][6] ;
 wire \core.cpuregs[18][7] ;
 wire \core.cpuregs[18][8] ;
 wire \core.cpuregs[18][9] ;
 wire \core.cpuregs[19][0] ;
 wire \core.cpuregs[19][10] ;
 wire \core.cpuregs[19][11] ;
 wire \core.cpuregs[19][12] ;
 wire \core.cpuregs[19][13] ;
 wire \core.cpuregs[19][14] ;
 wire \core.cpuregs[19][15] ;
 wire \core.cpuregs[19][16] ;
 wire \core.cpuregs[19][17] ;
 wire \core.cpuregs[19][18] ;
 wire \core.cpuregs[19][19] ;
 wire \core.cpuregs[19][1] ;
 wire \core.cpuregs[19][20] ;
 wire \core.cpuregs[19][21] ;
 wire \core.cpuregs[19][22] ;
 wire \core.cpuregs[19][23] ;
 wire \core.cpuregs[19][24] ;
 wire \core.cpuregs[19][25] ;
 wire \core.cpuregs[19][26] ;
 wire \core.cpuregs[19][27] ;
 wire \core.cpuregs[19][28] ;
 wire \core.cpuregs[19][29] ;
 wire \core.cpuregs[19][2] ;
 wire \core.cpuregs[19][30] ;
 wire \core.cpuregs[19][31] ;
 wire \core.cpuregs[19][3] ;
 wire \core.cpuregs[19][4] ;
 wire \core.cpuregs[19][5] ;
 wire \core.cpuregs[19][6] ;
 wire \core.cpuregs[19][7] ;
 wire \core.cpuregs[19][8] ;
 wire \core.cpuregs[19][9] ;
 wire \core.cpuregs[1][0] ;
 wire \core.cpuregs[1][10] ;
 wire \core.cpuregs[1][11] ;
 wire \core.cpuregs[1][12] ;
 wire \core.cpuregs[1][13] ;
 wire \core.cpuregs[1][14] ;
 wire \core.cpuregs[1][15] ;
 wire \core.cpuregs[1][16] ;
 wire \core.cpuregs[1][17] ;
 wire \core.cpuregs[1][18] ;
 wire \core.cpuregs[1][19] ;
 wire \core.cpuregs[1][1] ;
 wire \core.cpuregs[1][20] ;
 wire \core.cpuregs[1][21] ;
 wire \core.cpuregs[1][22] ;
 wire \core.cpuregs[1][23] ;
 wire \core.cpuregs[1][24] ;
 wire \core.cpuregs[1][25] ;
 wire \core.cpuregs[1][26] ;
 wire \core.cpuregs[1][27] ;
 wire \core.cpuregs[1][28] ;
 wire \core.cpuregs[1][29] ;
 wire \core.cpuregs[1][2] ;
 wire \core.cpuregs[1][30] ;
 wire \core.cpuregs[1][31] ;
 wire \core.cpuregs[1][3] ;
 wire \core.cpuregs[1][4] ;
 wire \core.cpuregs[1][5] ;
 wire \core.cpuregs[1][6] ;
 wire \core.cpuregs[1][7] ;
 wire \core.cpuregs[1][8] ;
 wire \core.cpuregs[1][9] ;
 wire \core.cpuregs[20][0] ;
 wire \core.cpuregs[20][10] ;
 wire \core.cpuregs[20][11] ;
 wire \core.cpuregs[20][12] ;
 wire \core.cpuregs[20][13] ;
 wire \core.cpuregs[20][14] ;
 wire \core.cpuregs[20][15] ;
 wire \core.cpuregs[20][16] ;
 wire \core.cpuregs[20][17] ;
 wire \core.cpuregs[20][18] ;
 wire \core.cpuregs[20][19] ;
 wire \core.cpuregs[20][1] ;
 wire \core.cpuregs[20][20] ;
 wire \core.cpuregs[20][21] ;
 wire \core.cpuregs[20][22] ;
 wire \core.cpuregs[20][23] ;
 wire \core.cpuregs[20][24] ;
 wire \core.cpuregs[20][25] ;
 wire \core.cpuregs[20][26] ;
 wire \core.cpuregs[20][27] ;
 wire \core.cpuregs[20][28] ;
 wire \core.cpuregs[20][29] ;
 wire \core.cpuregs[20][2] ;
 wire \core.cpuregs[20][30] ;
 wire \core.cpuregs[20][31] ;
 wire \core.cpuregs[20][3] ;
 wire \core.cpuregs[20][4] ;
 wire \core.cpuregs[20][5] ;
 wire \core.cpuregs[20][6] ;
 wire \core.cpuregs[20][7] ;
 wire \core.cpuregs[20][8] ;
 wire \core.cpuregs[20][9] ;
 wire \core.cpuregs[21][0] ;
 wire \core.cpuregs[21][10] ;
 wire \core.cpuregs[21][11] ;
 wire \core.cpuregs[21][12] ;
 wire \core.cpuregs[21][13] ;
 wire \core.cpuregs[21][14] ;
 wire \core.cpuregs[21][15] ;
 wire \core.cpuregs[21][16] ;
 wire \core.cpuregs[21][17] ;
 wire \core.cpuregs[21][18] ;
 wire \core.cpuregs[21][19] ;
 wire \core.cpuregs[21][1] ;
 wire \core.cpuregs[21][20] ;
 wire \core.cpuregs[21][21] ;
 wire \core.cpuregs[21][22] ;
 wire \core.cpuregs[21][23] ;
 wire \core.cpuregs[21][24] ;
 wire \core.cpuregs[21][25] ;
 wire \core.cpuregs[21][26] ;
 wire \core.cpuregs[21][27] ;
 wire \core.cpuregs[21][28] ;
 wire \core.cpuregs[21][29] ;
 wire \core.cpuregs[21][2] ;
 wire \core.cpuregs[21][30] ;
 wire \core.cpuregs[21][31] ;
 wire \core.cpuregs[21][3] ;
 wire \core.cpuregs[21][4] ;
 wire \core.cpuregs[21][5] ;
 wire \core.cpuregs[21][6] ;
 wire \core.cpuregs[21][7] ;
 wire \core.cpuregs[21][8] ;
 wire \core.cpuregs[21][9] ;
 wire \core.cpuregs[22][0] ;
 wire \core.cpuregs[22][10] ;
 wire \core.cpuregs[22][11] ;
 wire \core.cpuregs[22][12] ;
 wire \core.cpuregs[22][13] ;
 wire \core.cpuregs[22][14] ;
 wire \core.cpuregs[22][15] ;
 wire \core.cpuregs[22][16] ;
 wire \core.cpuregs[22][17] ;
 wire \core.cpuregs[22][18] ;
 wire \core.cpuregs[22][19] ;
 wire \core.cpuregs[22][1] ;
 wire \core.cpuregs[22][20] ;
 wire \core.cpuregs[22][21] ;
 wire \core.cpuregs[22][22] ;
 wire \core.cpuregs[22][23] ;
 wire \core.cpuregs[22][24] ;
 wire \core.cpuregs[22][25] ;
 wire \core.cpuregs[22][26] ;
 wire \core.cpuregs[22][27] ;
 wire \core.cpuregs[22][28] ;
 wire \core.cpuregs[22][29] ;
 wire \core.cpuregs[22][2] ;
 wire \core.cpuregs[22][30] ;
 wire \core.cpuregs[22][31] ;
 wire \core.cpuregs[22][3] ;
 wire \core.cpuregs[22][4] ;
 wire \core.cpuregs[22][5] ;
 wire \core.cpuregs[22][6] ;
 wire \core.cpuregs[22][7] ;
 wire \core.cpuregs[22][8] ;
 wire \core.cpuregs[22][9] ;
 wire \core.cpuregs[23][0] ;
 wire \core.cpuregs[23][10] ;
 wire \core.cpuregs[23][11] ;
 wire \core.cpuregs[23][12] ;
 wire \core.cpuregs[23][13] ;
 wire \core.cpuregs[23][14] ;
 wire \core.cpuregs[23][15] ;
 wire \core.cpuregs[23][16] ;
 wire \core.cpuregs[23][17] ;
 wire \core.cpuregs[23][18] ;
 wire \core.cpuregs[23][19] ;
 wire \core.cpuregs[23][1] ;
 wire \core.cpuregs[23][20] ;
 wire \core.cpuregs[23][21] ;
 wire \core.cpuregs[23][22] ;
 wire \core.cpuregs[23][23] ;
 wire \core.cpuregs[23][24] ;
 wire \core.cpuregs[23][25] ;
 wire \core.cpuregs[23][26] ;
 wire \core.cpuregs[23][27] ;
 wire \core.cpuregs[23][28] ;
 wire \core.cpuregs[23][29] ;
 wire \core.cpuregs[23][2] ;
 wire \core.cpuregs[23][30] ;
 wire \core.cpuregs[23][31] ;
 wire \core.cpuregs[23][3] ;
 wire \core.cpuregs[23][4] ;
 wire \core.cpuregs[23][5] ;
 wire \core.cpuregs[23][6] ;
 wire \core.cpuregs[23][7] ;
 wire \core.cpuregs[23][8] ;
 wire \core.cpuregs[23][9] ;
 wire \core.cpuregs[24][0] ;
 wire \core.cpuregs[24][10] ;
 wire \core.cpuregs[24][11] ;
 wire \core.cpuregs[24][12] ;
 wire \core.cpuregs[24][13] ;
 wire \core.cpuregs[24][14] ;
 wire \core.cpuregs[24][15] ;
 wire \core.cpuregs[24][16] ;
 wire \core.cpuregs[24][17] ;
 wire \core.cpuregs[24][18] ;
 wire \core.cpuregs[24][19] ;
 wire \core.cpuregs[24][1] ;
 wire \core.cpuregs[24][20] ;
 wire \core.cpuregs[24][21] ;
 wire \core.cpuregs[24][22] ;
 wire \core.cpuregs[24][23] ;
 wire \core.cpuregs[24][24] ;
 wire \core.cpuregs[24][25] ;
 wire \core.cpuregs[24][26] ;
 wire \core.cpuregs[24][27] ;
 wire \core.cpuregs[24][28] ;
 wire \core.cpuregs[24][29] ;
 wire \core.cpuregs[24][2] ;
 wire \core.cpuregs[24][30] ;
 wire \core.cpuregs[24][31] ;
 wire \core.cpuregs[24][3] ;
 wire \core.cpuregs[24][4] ;
 wire \core.cpuregs[24][5] ;
 wire \core.cpuregs[24][6] ;
 wire \core.cpuregs[24][7] ;
 wire \core.cpuregs[24][8] ;
 wire \core.cpuregs[24][9] ;
 wire \core.cpuregs[25][0] ;
 wire \core.cpuregs[25][10] ;
 wire \core.cpuregs[25][11] ;
 wire \core.cpuregs[25][12] ;
 wire \core.cpuregs[25][13] ;
 wire \core.cpuregs[25][14] ;
 wire \core.cpuregs[25][15] ;
 wire \core.cpuregs[25][16] ;
 wire \core.cpuregs[25][17] ;
 wire \core.cpuregs[25][18] ;
 wire \core.cpuregs[25][19] ;
 wire \core.cpuregs[25][1] ;
 wire \core.cpuregs[25][20] ;
 wire \core.cpuregs[25][21] ;
 wire \core.cpuregs[25][22] ;
 wire \core.cpuregs[25][23] ;
 wire \core.cpuregs[25][24] ;
 wire \core.cpuregs[25][25] ;
 wire \core.cpuregs[25][26] ;
 wire \core.cpuregs[25][27] ;
 wire \core.cpuregs[25][28] ;
 wire \core.cpuregs[25][29] ;
 wire \core.cpuregs[25][2] ;
 wire \core.cpuregs[25][30] ;
 wire \core.cpuregs[25][31] ;
 wire \core.cpuregs[25][3] ;
 wire \core.cpuregs[25][4] ;
 wire \core.cpuregs[25][5] ;
 wire \core.cpuregs[25][6] ;
 wire \core.cpuregs[25][7] ;
 wire \core.cpuregs[25][8] ;
 wire \core.cpuregs[25][9] ;
 wire \core.cpuregs[26][0] ;
 wire \core.cpuregs[26][10] ;
 wire \core.cpuregs[26][11] ;
 wire \core.cpuregs[26][12] ;
 wire \core.cpuregs[26][13] ;
 wire \core.cpuregs[26][14] ;
 wire \core.cpuregs[26][15] ;
 wire \core.cpuregs[26][16] ;
 wire \core.cpuregs[26][17] ;
 wire \core.cpuregs[26][18] ;
 wire \core.cpuregs[26][19] ;
 wire \core.cpuregs[26][1] ;
 wire \core.cpuregs[26][20] ;
 wire \core.cpuregs[26][21] ;
 wire \core.cpuregs[26][22] ;
 wire \core.cpuregs[26][23] ;
 wire \core.cpuregs[26][24] ;
 wire \core.cpuregs[26][25] ;
 wire \core.cpuregs[26][26] ;
 wire \core.cpuregs[26][27] ;
 wire \core.cpuregs[26][28] ;
 wire \core.cpuregs[26][29] ;
 wire \core.cpuregs[26][2] ;
 wire \core.cpuregs[26][30] ;
 wire \core.cpuregs[26][31] ;
 wire \core.cpuregs[26][3] ;
 wire \core.cpuregs[26][4] ;
 wire \core.cpuregs[26][5] ;
 wire \core.cpuregs[26][6] ;
 wire \core.cpuregs[26][7] ;
 wire \core.cpuregs[26][8] ;
 wire \core.cpuregs[26][9] ;
 wire \core.cpuregs[27][0] ;
 wire \core.cpuregs[27][10] ;
 wire \core.cpuregs[27][11] ;
 wire \core.cpuregs[27][12] ;
 wire \core.cpuregs[27][13] ;
 wire \core.cpuregs[27][14] ;
 wire \core.cpuregs[27][15] ;
 wire \core.cpuregs[27][16] ;
 wire \core.cpuregs[27][17] ;
 wire \core.cpuregs[27][18] ;
 wire \core.cpuregs[27][19] ;
 wire \core.cpuregs[27][1] ;
 wire \core.cpuregs[27][20] ;
 wire \core.cpuregs[27][21] ;
 wire \core.cpuregs[27][22] ;
 wire \core.cpuregs[27][23] ;
 wire \core.cpuregs[27][24] ;
 wire \core.cpuregs[27][25] ;
 wire \core.cpuregs[27][26] ;
 wire \core.cpuregs[27][27] ;
 wire \core.cpuregs[27][28] ;
 wire \core.cpuregs[27][29] ;
 wire \core.cpuregs[27][2] ;
 wire \core.cpuregs[27][30] ;
 wire \core.cpuregs[27][31] ;
 wire \core.cpuregs[27][3] ;
 wire \core.cpuregs[27][4] ;
 wire \core.cpuregs[27][5] ;
 wire \core.cpuregs[27][6] ;
 wire \core.cpuregs[27][7] ;
 wire \core.cpuregs[27][8] ;
 wire \core.cpuregs[27][9] ;
 wire \core.cpuregs[28][0] ;
 wire \core.cpuregs[28][10] ;
 wire \core.cpuregs[28][11] ;
 wire \core.cpuregs[28][12] ;
 wire \core.cpuregs[28][13] ;
 wire \core.cpuregs[28][14] ;
 wire \core.cpuregs[28][15] ;
 wire \core.cpuregs[28][16] ;
 wire \core.cpuregs[28][17] ;
 wire \core.cpuregs[28][18] ;
 wire \core.cpuregs[28][19] ;
 wire \core.cpuregs[28][1] ;
 wire \core.cpuregs[28][20] ;
 wire \core.cpuregs[28][21] ;
 wire \core.cpuregs[28][22] ;
 wire \core.cpuregs[28][23] ;
 wire \core.cpuregs[28][24] ;
 wire \core.cpuregs[28][25] ;
 wire \core.cpuregs[28][26] ;
 wire \core.cpuregs[28][27] ;
 wire \core.cpuregs[28][28] ;
 wire \core.cpuregs[28][29] ;
 wire \core.cpuregs[28][2] ;
 wire \core.cpuregs[28][30] ;
 wire \core.cpuregs[28][31] ;
 wire \core.cpuregs[28][3] ;
 wire \core.cpuregs[28][4] ;
 wire \core.cpuregs[28][5] ;
 wire \core.cpuregs[28][6] ;
 wire \core.cpuregs[28][7] ;
 wire \core.cpuregs[28][8] ;
 wire \core.cpuregs[28][9] ;
 wire \core.cpuregs[29][0] ;
 wire \core.cpuregs[29][10] ;
 wire \core.cpuregs[29][11] ;
 wire \core.cpuregs[29][12] ;
 wire \core.cpuregs[29][13] ;
 wire \core.cpuregs[29][14] ;
 wire \core.cpuregs[29][15] ;
 wire \core.cpuregs[29][16] ;
 wire \core.cpuregs[29][17] ;
 wire \core.cpuregs[29][18] ;
 wire \core.cpuregs[29][19] ;
 wire \core.cpuregs[29][1] ;
 wire \core.cpuregs[29][20] ;
 wire \core.cpuregs[29][21] ;
 wire \core.cpuregs[29][22] ;
 wire \core.cpuregs[29][23] ;
 wire \core.cpuregs[29][24] ;
 wire \core.cpuregs[29][25] ;
 wire \core.cpuregs[29][26] ;
 wire \core.cpuregs[29][27] ;
 wire \core.cpuregs[29][28] ;
 wire \core.cpuregs[29][29] ;
 wire \core.cpuregs[29][2] ;
 wire \core.cpuregs[29][30] ;
 wire \core.cpuregs[29][31] ;
 wire \core.cpuregs[29][3] ;
 wire \core.cpuregs[29][4] ;
 wire \core.cpuregs[29][5] ;
 wire \core.cpuregs[29][6] ;
 wire \core.cpuregs[29][7] ;
 wire \core.cpuregs[29][8] ;
 wire \core.cpuregs[29][9] ;
 wire \core.cpuregs[2][0] ;
 wire \core.cpuregs[2][10] ;
 wire \core.cpuregs[2][11] ;
 wire \core.cpuregs[2][12] ;
 wire \core.cpuregs[2][13] ;
 wire \core.cpuregs[2][14] ;
 wire \core.cpuregs[2][15] ;
 wire \core.cpuregs[2][16] ;
 wire \core.cpuregs[2][17] ;
 wire \core.cpuregs[2][18] ;
 wire \core.cpuregs[2][19] ;
 wire \core.cpuregs[2][1] ;
 wire \core.cpuregs[2][20] ;
 wire \core.cpuregs[2][21] ;
 wire \core.cpuregs[2][22] ;
 wire \core.cpuregs[2][23] ;
 wire \core.cpuregs[2][24] ;
 wire \core.cpuregs[2][25] ;
 wire \core.cpuregs[2][26] ;
 wire \core.cpuregs[2][27] ;
 wire \core.cpuregs[2][28] ;
 wire \core.cpuregs[2][29] ;
 wire \core.cpuregs[2][2] ;
 wire \core.cpuregs[2][30] ;
 wire \core.cpuregs[2][31] ;
 wire \core.cpuregs[2][3] ;
 wire \core.cpuregs[2][4] ;
 wire \core.cpuregs[2][5] ;
 wire \core.cpuregs[2][6] ;
 wire \core.cpuregs[2][7] ;
 wire \core.cpuregs[2][8] ;
 wire \core.cpuregs[2][9] ;
 wire \core.cpuregs[30][0] ;
 wire \core.cpuregs[30][10] ;
 wire \core.cpuregs[30][11] ;
 wire \core.cpuregs[30][12] ;
 wire \core.cpuregs[30][13] ;
 wire \core.cpuregs[30][14] ;
 wire \core.cpuregs[30][15] ;
 wire \core.cpuregs[30][16] ;
 wire \core.cpuregs[30][17] ;
 wire \core.cpuregs[30][18] ;
 wire \core.cpuregs[30][19] ;
 wire \core.cpuregs[30][1] ;
 wire \core.cpuregs[30][20] ;
 wire \core.cpuregs[30][21] ;
 wire \core.cpuregs[30][22] ;
 wire \core.cpuregs[30][23] ;
 wire \core.cpuregs[30][24] ;
 wire \core.cpuregs[30][25] ;
 wire \core.cpuregs[30][26] ;
 wire \core.cpuregs[30][27] ;
 wire \core.cpuregs[30][28] ;
 wire \core.cpuregs[30][29] ;
 wire \core.cpuregs[30][2] ;
 wire \core.cpuregs[30][30] ;
 wire \core.cpuregs[30][31] ;
 wire \core.cpuregs[30][3] ;
 wire \core.cpuregs[30][4] ;
 wire \core.cpuregs[30][5] ;
 wire \core.cpuregs[30][6] ;
 wire \core.cpuregs[30][7] ;
 wire \core.cpuregs[30][8] ;
 wire \core.cpuregs[30][9] ;
 wire \core.cpuregs[31][0] ;
 wire \core.cpuregs[31][10] ;
 wire \core.cpuregs[31][11] ;
 wire \core.cpuregs[31][12] ;
 wire \core.cpuregs[31][13] ;
 wire \core.cpuregs[31][14] ;
 wire \core.cpuregs[31][15] ;
 wire \core.cpuregs[31][16] ;
 wire \core.cpuregs[31][17] ;
 wire \core.cpuregs[31][18] ;
 wire \core.cpuregs[31][19] ;
 wire \core.cpuregs[31][1] ;
 wire \core.cpuregs[31][20] ;
 wire \core.cpuregs[31][21] ;
 wire \core.cpuregs[31][22] ;
 wire \core.cpuregs[31][23] ;
 wire \core.cpuregs[31][24] ;
 wire \core.cpuregs[31][25] ;
 wire \core.cpuregs[31][26] ;
 wire \core.cpuregs[31][27] ;
 wire \core.cpuregs[31][28] ;
 wire \core.cpuregs[31][29] ;
 wire \core.cpuregs[31][2] ;
 wire \core.cpuregs[31][30] ;
 wire \core.cpuregs[31][31] ;
 wire \core.cpuregs[31][3] ;
 wire \core.cpuregs[31][4] ;
 wire \core.cpuregs[31][5] ;
 wire \core.cpuregs[31][6] ;
 wire \core.cpuregs[31][7] ;
 wire \core.cpuregs[31][8] ;
 wire \core.cpuregs[31][9] ;
 wire \core.cpuregs[3][0] ;
 wire \core.cpuregs[3][10] ;
 wire \core.cpuregs[3][11] ;
 wire \core.cpuregs[3][12] ;
 wire \core.cpuregs[3][13] ;
 wire \core.cpuregs[3][14] ;
 wire \core.cpuregs[3][15] ;
 wire \core.cpuregs[3][16] ;
 wire \core.cpuregs[3][17] ;
 wire \core.cpuregs[3][18] ;
 wire \core.cpuregs[3][19] ;
 wire \core.cpuregs[3][1] ;
 wire \core.cpuregs[3][20] ;
 wire \core.cpuregs[3][21] ;
 wire \core.cpuregs[3][22] ;
 wire \core.cpuregs[3][23] ;
 wire \core.cpuregs[3][24] ;
 wire \core.cpuregs[3][25] ;
 wire \core.cpuregs[3][26] ;
 wire \core.cpuregs[3][27] ;
 wire \core.cpuregs[3][28] ;
 wire \core.cpuregs[3][29] ;
 wire \core.cpuregs[3][2] ;
 wire \core.cpuregs[3][30] ;
 wire \core.cpuregs[3][31] ;
 wire \core.cpuregs[3][3] ;
 wire \core.cpuregs[3][4] ;
 wire \core.cpuregs[3][5] ;
 wire \core.cpuregs[3][6] ;
 wire \core.cpuregs[3][7] ;
 wire \core.cpuregs[3][8] ;
 wire \core.cpuregs[3][9] ;
 wire \core.cpuregs[4][0] ;
 wire \core.cpuregs[4][10] ;
 wire \core.cpuregs[4][11] ;
 wire \core.cpuregs[4][12] ;
 wire \core.cpuregs[4][13] ;
 wire \core.cpuregs[4][14] ;
 wire \core.cpuregs[4][15] ;
 wire \core.cpuregs[4][16] ;
 wire \core.cpuregs[4][17] ;
 wire \core.cpuregs[4][18] ;
 wire \core.cpuregs[4][19] ;
 wire \core.cpuregs[4][1] ;
 wire \core.cpuregs[4][20] ;
 wire \core.cpuregs[4][21] ;
 wire \core.cpuregs[4][22] ;
 wire \core.cpuregs[4][23] ;
 wire \core.cpuregs[4][24] ;
 wire \core.cpuregs[4][25] ;
 wire \core.cpuregs[4][26] ;
 wire \core.cpuregs[4][27] ;
 wire \core.cpuregs[4][28] ;
 wire \core.cpuregs[4][29] ;
 wire \core.cpuregs[4][2] ;
 wire \core.cpuregs[4][30] ;
 wire \core.cpuregs[4][31] ;
 wire \core.cpuregs[4][3] ;
 wire \core.cpuregs[4][4] ;
 wire \core.cpuregs[4][5] ;
 wire \core.cpuregs[4][6] ;
 wire \core.cpuregs[4][7] ;
 wire \core.cpuregs[4][8] ;
 wire \core.cpuregs[4][9] ;
 wire \core.cpuregs[5][0] ;
 wire \core.cpuregs[5][10] ;
 wire \core.cpuregs[5][11] ;
 wire \core.cpuregs[5][12] ;
 wire \core.cpuregs[5][13] ;
 wire \core.cpuregs[5][14] ;
 wire \core.cpuregs[5][15] ;
 wire \core.cpuregs[5][16] ;
 wire \core.cpuregs[5][17] ;
 wire \core.cpuregs[5][18] ;
 wire \core.cpuregs[5][19] ;
 wire \core.cpuregs[5][1] ;
 wire \core.cpuregs[5][20] ;
 wire \core.cpuregs[5][21] ;
 wire \core.cpuregs[5][22] ;
 wire \core.cpuregs[5][23] ;
 wire \core.cpuregs[5][24] ;
 wire \core.cpuregs[5][25] ;
 wire \core.cpuregs[5][26] ;
 wire \core.cpuregs[5][27] ;
 wire \core.cpuregs[5][28] ;
 wire \core.cpuregs[5][29] ;
 wire \core.cpuregs[5][2] ;
 wire \core.cpuregs[5][30] ;
 wire \core.cpuregs[5][31] ;
 wire \core.cpuregs[5][3] ;
 wire \core.cpuregs[5][4] ;
 wire \core.cpuregs[5][5] ;
 wire \core.cpuregs[5][6] ;
 wire \core.cpuregs[5][7] ;
 wire \core.cpuregs[5][8] ;
 wire \core.cpuregs[5][9] ;
 wire \core.cpuregs[6][0] ;
 wire \core.cpuregs[6][10] ;
 wire \core.cpuregs[6][11] ;
 wire \core.cpuregs[6][12] ;
 wire \core.cpuregs[6][13] ;
 wire \core.cpuregs[6][14] ;
 wire \core.cpuregs[6][15] ;
 wire \core.cpuregs[6][16] ;
 wire \core.cpuregs[6][17] ;
 wire \core.cpuregs[6][18] ;
 wire \core.cpuregs[6][19] ;
 wire \core.cpuregs[6][1] ;
 wire \core.cpuregs[6][20] ;
 wire \core.cpuregs[6][21] ;
 wire \core.cpuregs[6][22] ;
 wire \core.cpuregs[6][23] ;
 wire \core.cpuregs[6][24] ;
 wire \core.cpuregs[6][25] ;
 wire \core.cpuregs[6][26] ;
 wire \core.cpuregs[6][27] ;
 wire \core.cpuregs[6][28] ;
 wire \core.cpuregs[6][29] ;
 wire \core.cpuregs[6][2] ;
 wire \core.cpuregs[6][30] ;
 wire \core.cpuregs[6][31] ;
 wire \core.cpuregs[6][3] ;
 wire \core.cpuregs[6][4] ;
 wire \core.cpuregs[6][5] ;
 wire \core.cpuregs[6][6] ;
 wire \core.cpuregs[6][7] ;
 wire \core.cpuregs[6][8] ;
 wire \core.cpuregs[6][9] ;
 wire \core.cpuregs[7][0] ;
 wire \core.cpuregs[7][10] ;
 wire \core.cpuregs[7][11] ;
 wire \core.cpuregs[7][12] ;
 wire \core.cpuregs[7][13] ;
 wire \core.cpuregs[7][14] ;
 wire \core.cpuregs[7][15] ;
 wire \core.cpuregs[7][16] ;
 wire \core.cpuregs[7][17] ;
 wire \core.cpuregs[7][18] ;
 wire \core.cpuregs[7][19] ;
 wire \core.cpuregs[7][1] ;
 wire \core.cpuregs[7][20] ;
 wire \core.cpuregs[7][21] ;
 wire \core.cpuregs[7][22] ;
 wire \core.cpuregs[7][23] ;
 wire \core.cpuregs[7][24] ;
 wire \core.cpuregs[7][25] ;
 wire \core.cpuregs[7][26] ;
 wire \core.cpuregs[7][27] ;
 wire \core.cpuregs[7][28] ;
 wire \core.cpuregs[7][29] ;
 wire \core.cpuregs[7][2] ;
 wire \core.cpuregs[7][30] ;
 wire \core.cpuregs[7][31] ;
 wire \core.cpuregs[7][3] ;
 wire \core.cpuregs[7][4] ;
 wire \core.cpuregs[7][5] ;
 wire \core.cpuregs[7][6] ;
 wire \core.cpuregs[7][7] ;
 wire \core.cpuregs[7][8] ;
 wire \core.cpuregs[7][9] ;
 wire \core.cpuregs[8][0] ;
 wire \core.cpuregs[8][10] ;
 wire \core.cpuregs[8][11] ;
 wire \core.cpuregs[8][12] ;
 wire \core.cpuregs[8][13] ;
 wire \core.cpuregs[8][14] ;
 wire \core.cpuregs[8][15] ;
 wire \core.cpuregs[8][16] ;
 wire \core.cpuregs[8][17] ;
 wire \core.cpuregs[8][18] ;
 wire \core.cpuregs[8][19] ;
 wire \core.cpuregs[8][1] ;
 wire \core.cpuregs[8][20] ;
 wire \core.cpuregs[8][21] ;
 wire \core.cpuregs[8][22] ;
 wire \core.cpuregs[8][23] ;
 wire \core.cpuregs[8][24] ;
 wire \core.cpuregs[8][25] ;
 wire \core.cpuregs[8][26] ;
 wire \core.cpuregs[8][27] ;
 wire \core.cpuregs[8][28] ;
 wire \core.cpuregs[8][29] ;
 wire \core.cpuregs[8][2] ;
 wire \core.cpuregs[8][30] ;
 wire \core.cpuregs[8][31] ;
 wire \core.cpuregs[8][3] ;
 wire \core.cpuregs[8][4] ;
 wire \core.cpuregs[8][5] ;
 wire \core.cpuregs[8][6] ;
 wire \core.cpuregs[8][7] ;
 wire \core.cpuregs[8][8] ;
 wire \core.cpuregs[8][9] ;
 wire \core.cpuregs[9][0] ;
 wire \core.cpuregs[9][10] ;
 wire \core.cpuregs[9][11] ;
 wire \core.cpuregs[9][12] ;
 wire \core.cpuregs[9][13] ;
 wire \core.cpuregs[9][14] ;
 wire \core.cpuregs[9][15] ;
 wire \core.cpuregs[9][16] ;
 wire \core.cpuregs[9][17] ;
 wire \core.cpuregs[9][18] ;
 wire \core.cpuregs[9][19] ;
 wire \core.cpuregs[9][1] ;
 wire \core.cpuregs[9][20] ;
 wire \core.cpuregs[9][21] ;
 wire \core.cpuregs[9][22] ;
 wire \core.cpuregs[9][23] ;
 wire \core.cpuregs[9][24] ;
 wire \core.cpuregs[9][25] ;
 wire \core.cpuregs[9][26] ;
 wire \core.cpuregs[9][27] ;
 wire \core.cpuregs[9][28] ;
 wire \core.cpuregs[9][29] ;
 wire \core.cpuregs[9][2] ;
 wire \core.cpuregs[9][30] ;
 wire \core.cpuregs[9][31] ;
 wire \core.cpuregs[9][3] ;
 wire \core.cpuregs[9][4] ;
 wire \core.cpuregs[9][5] ;
 wire \core.cpuregs[9][6] ;
 wire \core.cpuregs[9][7] ;
 wire \core.cpuregs[9][8] ;
 wire \core.cpuregs[9][9] ;
 wire \core.decoded_imm[0] ;
 wire \core.decoded_imm[10] ;
 wire \core.decoded_imm[11] ;
 wire \core.decoded_imm[12] ;
 wire \core.decoded_imm[13] ;
 wire \core.decoded_imm[14] ;
 wire \core.decoded_imm[15] ;
 wire \core.decoded_imm[16] ;
 wire \core.decoded_imm[17] ;
 wire \core.decoded_imm[18] ;
 wire \core.decoded_imm[19] ;
 wire \core.decoded_imm[1] ;
 wire \core.decoded_imm[20] ;
 wire \core.decoded_imm[21] ;
 wire \core.decoded_imm[22] ;
 wire \core.decoded_imm[23] ;
 wire \core.decoded_imm[24] ;
 wire \core.decoded_imm[25] ;
 wire \core.decoded_imm[26] ;
 wire \core.decoded_imm[27] ;
 wire \core.decoded_imm[28] ;
 wire \core.decoded_imm[29] ;
 wire \core.decoded_imm[2] ;
 wire \core.decoded_imm[30] ;
 wire \core.decoded_imm[31] ;
 wire \core.decoded_imm[3] ;
 wire \core.decoded_imm[4] ;
 wire \core.decoded_imm[5] ;
 wire \core.decoded_imm[6] ;
 wire \core.decoded_imm[7] ;
 wire \core.decoded_imm[8] ;
 wire \core.decoded_imm[9] ;
 wire \core.decoded_imm_j[10] ;
 wire \core.decoded_imm_j[11] ;
 wire \core.decoded_imm_j[12] ;
 wire \core.decoded_imm_j[13] ;
 wire \core.decoded_imm_j[14] ;
 wire \core.decoded_imm_j[15] ;
 wire \core.decoded_imm_j[16] ;
 wire \core.decoded_imm_j[17] ;
 wire \core.decoded_imm_j[18] ;
 wire \core.decoded_imm_j[19] ;
 wire \core.decoded_imm_j[1] ;
 wire \core.decoded_imm_j[20] ;
 wire \core.decoded_imm_j[2] ;
 wire \core.decoded_imm_j[3] ;
 wire \core.decoded_imm_j[4] ;
 wire \core.decoded_imm_j[5] ;
 wire \core.decoded_imm_j[6] ;
 wire \core.decoded_imm_j[7] ;
 wire \core.decoded_imm_j[8] ;
 wire \core.decoded_imm_j[9] ;
 wire \core.decoded_rd[0] ;
 wire \core.decoded_rd[1] ;
 wire \core.decoded_rd[2] ;
 wire \core.decoded_rd[3] ;
 wire \core.decoded_rd[4] ;
 wire \core.decoder_pseudo_trigger ;
 wire \core.decoder_trigger ;
 wire \core.instr_add ;
 wire \core.instr_addi ;
 wire \core.instr_and ;
 wire \core.instr_andi ;
 wire \core.instr_auipc ;
 wire \core.instr_beq ;
 wire \core.instr_bge ;
 wire \core.instr_bgeu ;
 wire \core.instr_blt ;
 wire \core.instr_bltu ;
 wire \core.instr_bne ;
 wire \core.instr_fence ;
 wire \core.instr_jal ;
 wire \core.instr_jalr ;
 wire \core.instr_lb ;
 wire \core.instr_lbu ;
 wire \core.instr_lh ;
 wire \core.instr_lhu ;
 wire \core.instr_lui ;
 wire \core.instr_lw ;
 wire \core.instr_or ;
 wire \core.instr_ori ;
 wire \core.instr_rdcycle ;
 wire \core.instr_rdcycleh ;
 wire \core.instr_rdinstr ;
 wire \core.instr_rdinstrh ;
 wire \core.instr_sb ;
 wire \core.instr_sh ;
 wire \core.instr_sll ;
 wire \core.instr_slli ;
 wire \core.instr_slt ;
 wire \core.instr_slti ;
 wire \core.instr_sltiu ;
 wire \core.instr_sltu ;
 wire \core.instr_sra ;
 wire \core.instr_srai ;
 wire \core.instr_srl ;
 wire \core.instr_srli ;
 wire \core.instr_sub ;
 wire \core.instr_sw ;
 wire \core.instr_xor ;
 wire \core.instr_xori ;
 wire \core.is_alu_reg_imm ;
 wire \core.is_alu_reg_reg ;
 wire \core.is_beq_bne_blt_bge_bltu_bgeu ;
 wire \core.is_compare ;
 wire \core.is_jalr_addi_slti_sltiu_xori_ori_andi ;
 wire \core.is_lb_lh_lw_lbu_lhu ;
 wire \core.is_lui_auipc_jal ;
 wire \core.is_sb_sh_sw ;
 wire \core.is_sll_srl_sra ;
 wire \core.is_slli_srli_srai ;
 wire \core.is_slti_blt_slt ;
 wire \core.is_sltiu_bltu_sltu ;
 wire \core.latched_branch ;
 wire \core.latched_is_lb ;
 wire \core.latched_is_lh ;
 wire \core.latched_rd[0] ;
 wire \core.latched_rd[1] ;
 wire \core.latched_rd[2] ;
 wire \core.latched_rd[3] ;
 wire \core.latched_rd[4] ;
 wire \core.latched_stalu ;
 wire \core.latched_store ;
 wire \core.mem_do_prefetch ;
 wire \core.mem_do_rdata ;
 wire \core.mem_do_rinst ;
 wire \core.mem_do_wdata ;
 wire \core.mem_la_wdata[0] ;
 wire \core.mem_la_wdata[1] ;
 wire \core.mem_la_wdata[2] ;
 wire \core.mem_la_wdata[3] ;
 wire \core.mem_la_wdata[4] ;
 wire \core.mem_la_wdata[5] ;
 wire \core.mem_la_wdata[6] ;
 wire \core.mem_la_wdata[7] ;
 wire \core.mem_rdata_q[0] ;
 wire \core.mem_rdata_q[10] ;
 wire \core.mem_rdata_q[11] ;
 wire \core.mem_rdata_q[12] ;
 wire \core.mem_rdata_q[13] ;
 wire \core.mem_rdata_q[14] ;
 wire \core.mem_rdata_q[15] ;
 wire \core.mem_rdata_q[16] ;
 wire \core.mem_rdata_q[17] ;
 wire \core.mem_rdata_q[18] ;
 wire \core.mem_rdata_q[19] ;
 wire \core.mem_rdata_q[1] ;
 wire \core.mem_rdata_q[20] ;
 wire \core.mem_rdata_q[21] ;
 wire \core.mem_rdata_q[22] ;
 wire \core.mem_rdata_q[23] ;
 wire \core.mem_rdata_q[24] ;
 wire \core.mem_rdata_q[25] ;
 wire \core.mem_rdata_q[26] ;
 wire \core.mem_rdata_q[27] ;
 wire \core.mem_rdata_q[28] ;
 wire \core.mem_rdata_q[29] ;
 wire \core.mem_rdata_q[2] ;
 wire \core.mem_rdata_q[30] ;
 wire \core.mem_rdata_q[31] ;
 wire \core.mem_rdata_q[3] ;
 wire \core.mem_rdata_q[4] ;
 wire \core.mem_rdata_q[5] ;
 wire \core.mem_rdata_q[6] ;
 wire \core.mem_rdata_q[7] ;
 wire \core.mem_rdata_q[8] ;
 wire \core.mem_rdata_q[9] ;
 wire \core.mem_state[0] ;
 wire \core.mem_state[1] ;
 wire \core.mem_wordsize[0] ;
 wire \core.mem_wordsize[1] ;
 wire \core.mem_wordsize[2] ;
 wire \core.pcpi_rs1[0] ;
 wire \core.pcpi_rs1[10] ;
 wire \core.pcpi_rs1[11] ;
 wire \core.pcpi_rs1[12] ;
 wire \core.pcpi_rs1[13] ;
 wire \core.pcpi_rs1[14] ;
 wire \core.pcpi_rs1[15] ;
 wire \core.pcpi_rs1[16] ;
 wire \core.pcpi_rs1[17] ;
 wire \core.pcpi_rs1[18] ;
 wire \core.pcpi_rs1[19] ;
 wire \core.pcpi_rs1[1] ;
 wire \core.pcpi_rs1[20] ;
 wire \core.pcpi_rs1[21] ;
 wire \core.pcpi_rs1[22] ;
 wire \core.pcpi_rs1[23] ;
 wire \core.pcpi_rs1[24] ;
 wire \core.pcpi_rs1[25] ;
 wire \core.pcpi_rs1[26] ;
 wire \core.pcpi_rs1[27] ;
 wire \core.pcpi_rs1[28] ;
 wire \core.pcpi_rs1[29] ;
 wire \core.pcpi_rs1[2] ;
 wire \core.pcpi_rs1[30] ;
 wire \core.pcpi_rs1[31] ;
 wire \core.pcpi_rs1[3] ;
 wire \core.pcpi_rs1[4] ;
 wire \core.pcpi_rs1[5] ;
 wire \core.pcpi_rs1[6] ;
 wire \core.pcpi_rs1[7] ;
 wire \core.pcpi_rs1[8] ;
 wire \core.pcpi_rs1[9] ;
 wire \core.pcpi_rs2[10] ;
 wire \core.pcpi_rs2[11] ;
 wire \core.pcpi_rs2[12] ;
 wire \core.pcpi_rs2[13] ;
 wire \core.pcpi_rs2[14] ;
 wire \core.pcpi_rs2[15] ;
 wire \core.pcpi_rs2[16] ;
 wire \core.pcpi_rs2[17] ;
 wire \core.pcpi_rs2[18] ;
 wire \core.pcpi_rs2[19] ;
 wire \core.pcpi_rs2[20] ;
 wire \core.pcpi_rs2[21] ;
 wire \core.pcpi_rs2[22] ;
 wire \core.pcpi_rs2[23] ;
 wire \core.pcpi_rs2[24] ;
 wire \core.pcpi_rs2[25] ;
 wire \core.pcpi_rs2[26] ;
 wire \core.pcpi_rs2[27] ;
 wire \core.pcpi_rs2[28] ;
 wire \core.pcpi_rs2[29] ;
 wire \core.pcpi_rs2[30] ;
 wire \core.pcpi_rs2[31] ;
 wire \core.pcpi_rs2[8] ;
 wire \core.pcpi_rs2[9] ;
 wire \core.reg_next_pc[10] ;
 wire \core.reg_next_pc[11] ;
 wire \core.reg_next_pc[12] ;
 wire \core.reg_next_pc[13] ;
 wire \core.reg_next_pc[14] ;
 wire \core.reg_next_pc[15] ;
 wire \core.reg_next_pc[16] ;
 wire \core.reg_next_pc[17] ;
 wire \core.reg_next_pc[18] ;
 wire \core.reg_next_pc[19] ;
 wire \core.reg_next_pc[1] ;
 wire \core.reg_next_pc[20] ;
 wire \core.reg_next_pc[21] ;
 wire \core.reg_next_pc[22] ;
 wire \core.reg_next_pc[23] ;
 wire \core.reg_next_pc[24] ;
 wire \core.reg_next_pc[25] ;
 wire \core.reg_next_pc[26] ;
 wire \core.reg_next_pc[27] ;
 wire \core.reg_next_pc[28] ;
 wire \core.reg_next_pc[29] ;
 wire \core.reg_next_pc[2] ;
 wire \core.reg_next_pc[30] ;
 wire \core.reg_next_pc[31] ;
 wire \core.reg_next_pc[3] ;
 wire \core.reg_next_pc[4] ;
 wire \core.reg_next_pc[5] ;
 wire \core.reg_next_pc[6] ;
 wire \core.reg_next_pc[7] ;
 wire \core.reg_next_pc[8] ;
 wire \core.reg_next_pc[9] ;
 wire \core.reg_out[0] ;
 wire \core.reg_out[10] ;
 wire \core.reg_out[11] ;
 wire \core.reg_out[12] ;
 wire \core.reg_out[13] ;
 wire \core.reg_out[14] ;
 wire \core.reg_out[15] ;
 wire \core.reg_out[16] ;
 wire \core.reg_out[17] ;
 wire \core.reg_out[18] ;
 wire \core.reg_out[19] ;
 wire \core.reg_out[1] ;
 wire \core.reg_out[20] ;
 wire \core.reg_out[21] ;
 wire \core.reg_out[22] ;
 wire \core.reg_out[23] ;
 wire \core.reg_out[24] ;
 wire \core.reg_out[25] ;
 wire \core.reg_out[26] ;
 wire \core.reg_out[27] ;
 wire \core.reg_out[28] ;
 wire \core.reg_out[29] ;
 wire \core.reg_out[2] ;
 wire \core.reg_out[30] ;
 wire \core.reg_out[31] ;
 wire \core.reg_out[3] ;
 wire \core.reg_out[4] ;
 wire \core.reg_out[5] ;
 wire \core.reg_out[6] ;
 wire \core.reg_out[7] ;
 wire \core.reg_out[8] ;
 wire \core.reg_out[9] ;
 wire \core.reg_pc[10] ;
 wire \core.reg_pc[11] ;
 wire \core.reg_pc[12] ;
 wire \core.reg_pc[13] ;
 wire \core.reg_pc[14] ;
 wire \core.reg_pc[15] ;
 wire \core.reg_pc[16] ;
 wire \core.reg_pc[17] ;
 wire \core.reg_pc[18] ;
 wire \core.reg_pc[19] ;
 wire \core.reg_pc[1] ;
 wire \core.reg_pc[20] ;
 wire \core.reg_pc[21] ;
 wire \core.reg_pc[22] ;
 wire \core.reg_pc[23] ;
 wire \core.reg_pc[24] ;
 wire \core.reg_pc[25] ;
 wire \core.reg_pc[26] ;
 wire \core.reg_pc[27] ;
 wire \core.reg_pc[28] ;
 wire \core.reg_pc[29] ;
 wire \core.reg_pc[2] ;
 wire \core.reg_pc[30] ;
 wire \core.reg_pc[31] ;
 wire \core.reg_pc[3] ;
 wire \core.reg_pc[4] ;
 wire \core.reg_pc[5] ;
 wire \core.reg_pc[6] ;
 wire \core.reg_pc[7] ;
 wire \core.reg_pc[8] ;
 wire \core.reg_pc[9] ;
 wire \core.reg_sh[0] ;
 wire \core.reg_sh[1] ;
 wire \core.reg_sh[2] ;
 wire \core.reg_sh[3] ;
 wire \core.reg_sh[4] ;

 sky130_fd_sc_hd__or3_2 _07548_ (.A(\core.instr_sltu ),
    .B(\core.instr_bltu ),
    .C(\core.instr_sltiu ),
    .X(_02016_));
 sky130_fd_sc_hd__buf_1 _07549_ (.A(_02016_),
    .X(_00033_));
 sky130_fd_sc_hd__or3_2 _07550_ (.A(\core.instr_slt ),
    .B(\core.instr_blt ),
    .C(\core.instr_slti ),
    .X(_02017_));
 sky130_fd_sc_hd__buf_1 _07551_ (.A(_02017_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_1 _07552_ (.A(\core.instr_jal ),
    .X(_02018_));
 sky130_fd_sc_hd__buf_1 _07553_ (.A(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__or2_2 _07554_ (.A(\core.instr_auipc ),
    .B(\core.instr_lui ),
    .X(_02020_));
 sky130_fd_sc_hd__buf_1 _07555_ (.A(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__or2_2 _07556_ (.A(_02019_),
    .B(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__buf_1 _07557_ (.A(_02022_),
    .X(_00031_));
 sky130_fd_sc_hd__buf_1 _07558_ (.A(\core.mem_wordsize[1] ),
    .X(_02023_));
 sky130_fd_sc_hd__buf_1 _07559_ (.A(resetn),
    .X(_02024_));
 sky130_fd_sc_hd__and2_2 _07560_ (.A(mem_valid),
    .B(mem_ready),
    .X(_02025_));
 sky130_fd_sc_hd__buf_1 _07561_ (.A(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__or2_2 _07562_ (.A(\core.mem_state[1] ),
    .B(\core.mem_state[0] ),
    .X(_02027_));
 sky130_fd_sc_hd__o311a_2 _07563_ (.A1(\core.mem_do_rinst ),
    .A2(\core.mem_do_rdata ),
    .A3(\core.mem_do_wdata ),
    .B1(_02026_),
    .C1(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__a31o_2 _07564_ (.A1(\core.mem_do_rinst ),
    .A2(\core.mem_state[1] ),
    .A3(\core.mem_state[0] ),
    .B1(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_2 _07565_ (.A(_02024_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__and2_2 _07566_ (.A(\core.mem_do_prefetch ),
    .B(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__nor2_2 _07567_ (.A(\core.mem_do_wdata ),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_2 _07568_ (.A(\core.cpu_state[5] ),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__or3_2 _07569_ (.A(\core.instr_sb ),
    .B(\core.instr_sw ),
    .C(\core.instr_sh ),
    .X(_02034_));
 sky130_fd_sc_hd__or2_2 _07570_ (.A(_02033_),
    .B(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__inv_2 _07571_ (.A(\core.cpu_state[6] ),
    .Y(_02036_));
 sky130_fd_sc_hd__or2_2 _07572_ (.A(\core.mem_do_rdata ),
    .B(_02031_),
    .X(_02037_));
 sky130_fd_sc_hd__or4_2 _07573_ (.A(\core.instr_lb ),
    .B(\core.instr_lbu ),
    .C(\core.instr_lh ),
    .D(\core.instr_lhu ),
    .X(_02038_));
 sky130_fd_sc_hd__or4_2 _07574_ (.A(_02036_),
    .B(\core.instr_lw ),
    .C(_02037_),
    .D(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__or2_2 _07575_ (.A(\core.cpu_state[6] ),
    .B(\core.cpu_state[5] ),
    .X(_02040_));
 sky130_fd_sc_hd__buf_1 _07576_ (.A(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__buf_1 _07577_ (.A(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__o21ai_2 _07578_ (.A1(\core.mem_do_wdata ),
    .A2(_02031_),
    .B1(\core.cpu_state[5] ),
    .Y(_02043_));
 sky130_fd_sc_hd__o211a_2 _07579_ (.A1(\core.cpu_state[1] ),
    .A2(_02042_),
    .B1(_02043_),
    .C1(_02024_),
    .X(_02044_));
 sky130_fd_sc_hd__buf_1 _07580_ (.A(\core.cpu_state[6] ),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_2 _07581_ (.A(_02045_),
    .B(_02037_),
    .Y(_02046_));
 sky130_fd_sc_hd__nand4_2 _07582_ (.A(_02035_),
    .B(_02039_),
    .C(_02044_),
    .D(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__inv_2 _07583_ (.A(resetn),
    .Y(_02048_));
 sky130_fd_sc_hd__buf_1 _07584_ (.A(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__nor2_2 _07585_ (.A(_02049_),
    .B(_02033_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor2_2 _07586_ (.A(_02036_),
    .B(_02037_),
    .Y(_02051_));
 sky130_fd_sc_hd__buf_1 _07587_ (.A(_02024_),
    .X(_02052_));
 sky130_fd_sc_hd__o211a_2 _07588_ (.A1(\core.instr_lb ),
    .A2(\core.instr_lbu ),
    .B1(_02051_),
    .C1(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__a221o_2 _07589_ (.A1(_02023_),
    .A2(_02047_),
    .B1(_02050_),
    .B2(\core.instr_sb ),
    .C1(_02053_),
    .X(_00018_));
 sky130_fd_sc_hd__buf_1 _07590_ (.A(_02048_),
    .X(_02054_));
 sky130_fd_sc_hd__buf_1 _07591_ (.A(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__inv_2 _07592_ (.A(\core.cpu_state[2] ),
    .Y(_02056_));
 sky130_fd_sc_hd__or4_2 _07593_ (.A(\core.instr_rdinstr ),
    .B(\core.instr_rdinstrh ),
    .C(\core.instr_rdcycle ),
    .D(\core.instr_rdcycleh ),
    .X(_02057_));
 sky130_fd_sc_hd__or2_2 _07594_ (.A(\core.instr_bgeu ),
    .B(\core.instr_bge ),
    .X(_02058_));
 sky130_fd_sc_hd__or2_2 _07595_ (.A(\core.instr_sra ),
    .B(\core.instr_srai ),
    .X(_02059_));
 sky130_fd_sc_hd__or4_2 _07596_ (.A(\core.instr_sll ),
    .B(\core.instr_slli ),
    .C(_02058_),
    .D(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__or4_2 _07597_ (.A(\core.instr_andi ),
    .B(\core.instr_sub ),
    .C(\core.instr_srl ),
    .D(\core.instr_or ),
    .X(_02061_));
 sky130_fd_sc_hd__or4_2 _07598_ (.A(\core.instr_addi ),
    .B(\core.instr_xori ),
    .C(_02020_),
    .D(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__or3_2 _07599_ (.A(\core.instr_jal ),
    .B(\core.instr_jalr ),
    .C(\core.instr_lw ),
    .X(_02063_));
 sky130_fd_sc_hd__or4_2 _07600_ (.A(\core.instr_ori ),
    .B(\core.instr_beq ),
    .C(\core.instr_bne ),
    .D(\core.instr_srli ),
    .X(_02064_));
 sky130_fd_sc_hd__or4_2 _07601_ (.A(\core.instr_and ),
    .B(\core.instr_fence ),
    .C(\core.instr_xor ),
    .D(\core.instr_add ),
    .X(_02065_));
 sky130_fd_sc_hd__or4_2 _07602_ (.A(_00033_),
    .B(_02063_),
    .C(_02064_),
    .D(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__or4_2 _07603_ (.A(_00032_),
    .B(_02034_),
    .C(_02038_),
    .D(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__or4_2 _07604_ (.A(_02057_),
    .B(_02060_),
    .C(_02062_),
    .D(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__buf_1 _07605_ (.A(\core.mem_wordsize[2] ),
    .X(_02069_));
 sky130_fd_sc_hd__buf_1 _07606_ (.A(\core.pcpi_rs1[0] ),
    .X(_02070_));
 sky130_fd_sc_hd__buf_1 _07607_ (.A(\core.pcpi_rs1[1] ),
    .X(_02071_));
 sky130_fd_sc_hd__or2_2 _07608_ (.A(_02070_),
    .B(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a22o_2 _07609_ (.A1(_02069_),
    .A2(_02070_),
    .B1(\core.mem_wordsize[0] ),
    .B2(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__o21a_2 _07610_ (.A1(\core.mem_do_rdata ),
    .A2(\core.mem_do_wdata ),
    .B1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__a21oi_2 _07611_ (.A1(\core.mem_do_rinst ),
    .A2(\core.reg_pc[1] ),
    .B1(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__inv_2 _07612_ (.A(\core.cpu_state[0] ),
    .Y(_02076_));
 sky130_fd_sc_hd__o211a_2 _07613_ (.A1(_02056_),
    .A2(_02068_),
    .B1(_02075_),
    .C1(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__nor2_2 _07614_ (.A(_02055_),
    .B(_02077_),
    .Y(_00010_));
 sky130_fd_sc_hd__and3_2 _07615_ (.A(\core.cpu_state[5] ),
    .B(\core.instr_sw ),
    .C(_02032_),
    .X(_02078_));
 sky130_fd_sc_hd__buf_1 _07616_ (.A(\core.cpu_state[1] ),
    .X(_02079_));
 sky130_fd_sc_hd__buf_1 _07617_ (.A(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__a211o_2 _07618_ (.A1(\core.instr_lw ),
    .A2(_02051_),
    .B1(_02078_),
    .C1(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__buf_1 _07619_ (.A(_02052_),
    .X(_02082_));
 sky130_fd_sc_hd__buf_1 _07620_ (.A(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a22o_2 _07621_ (.A1(\core.mem_wordsize[0] ),
    .A2(_02047_),
    .B1(_02081_),
    .B2(_02083_),
    .X(_00017_));
 sky130_fd_sc_hd__and2_2 _07622_ (.A(_02024_),
    .B(_02075_),
    .X(_02084_));
 sky130_fd_sc_hd__and2_2 _07623_ (.A(\core.is_lb_lh_lw_lbu_lhu ),
    .B(_02068_),
    .X(_02085_));
 sky130_fd_sc_hd__or2_2 _07624_ (.A(\core.mem_do_prefetch ),
    .B(_02030_),
    .X(_02086_));
 sky130_fd_sc_hd__buf_1 _07625_ (.A(_02045_),
    .X(_02087_));
 sky130_fd_sc_hd__a22o_2 _07626_ (.A1(\core.cpu_state[2] ),
    .A2(_02085_),
    .B1(_02086_),
    .B2(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__and2_2 _07627_ (.A(_02084_),
    .B(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__buf_1 _07628_ (.A(_02089_),
    .X(_00016_));
 sky130_fd_sc_hd__buf_1 _07629_ (.A(\core.is_sb_sh_sw ),
    .X(_02090_));
 sky130_fd_sc_hd__buf_1 _07630_ (.A(\core.is_lb_lh_lw_lbu_lhu ),
    .X(_02091_));
 sky130_fd_sc_hd__or3b_2 _07631_ (.A(\core.is_slli_srli_srai ),
    .B(_02057_),
    .C_N(_02068_),
    .X(_02092_));
 sky130_fd_sc_hd__nor3_2 _07632_ (.A(_02056_),
    .B(_02091_),
    .C(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_2 _07633_ (.A(\core.is_lui_auipc_jal ),
    .B(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .Y(_02094_));
 sky130_fd_sc_hd__buf_1 _07634_ (.A(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__a32o_2 _07635_ (.A1(_02090_),
    .A2(_02093_),
    .A3(_02095_),
    .B1(_02086_),
    .B2(\core.cpu_state[5] ),
    .X(_02096_));
 sky130_fd_sc_hd__and2_2 _07636_ (.A(_02084_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__buf_1 _07637_ (.A(_02097_),
    .X(_00015_));
 sky130_fd_sc_hd__or3_2 _07638_ (.A(\core.reg_sh[4] ),
    .B(\core.reg_sh[3] ),
    .C(\core.reg_sh[2] ),
    .X(_02098_));
 sky130_fd_sc_hd__buf_1 _07639_ (.A(_02098_),
    .X(_02099_));
 sky130_fd_sc_hd__or3_2 _07640_ (.A(\core.reg_sh[0] ),
    .B(\core.reg_sh[1] ),
    .C(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__nand2_2 _07641_ (.A(\core.cpu_state[4] ),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__inv_2 _07642_ (.A(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__a32o_2 _07643_ (.A1(\core.is_sll_srl_sra ),
    .A2(_02093_),
    .A3(_02095_),
    .B1(\core.is_slli_srli_srai ),
    .B2(\core.cpu_state[2] ),
    .X(_02103_));
 sky130_fd_sc_hd__o21a_2 _07644_ (.A1(_02102_),
    .A2(_02103_),
    .B1(_02084_),
    .X(_00014_));
 sky130_fd_sc_hd__or4_2 _07645_ (.A(_02090_),
    .B(_02091_),
    .C(\core.is_sll_srl_sra ),
    .D(_02092_),
    .X(_02104_));
 sky130_fd_sc_hd__nand2_2 _07646_ (.A(_02095_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__a32o_2 _07647_ (.A1(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(\core.cpu_state[3] ),
    .A3(_02030_),
    .B1(_02105_),
    .B2(\core.cpu_state[2] ),
    .X(_02106_));
 sky130_fd_sc_hd__and2_2 _07648_ (.A(_02084_),
    .B(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__buf_1 _07649_ (.A(_02107_),
    .X(_00013_));
 sky130_fd_sc_hd__inv_2 _07650_ (.A(\core.decoder_trigger ),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_2 _07651_ (.A(_02108_),
    .B(\core.instr_jal ),
    .Y(_02109_));
 sky130_fd_sc_hd__inv_2 _07652_ (.A(\core.cpu_state[1] ),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_2 _07653_ (.A(_02110_),
    .B(_02048_),
    .Y(_02111_));
 sky130_fd_sc_hd__and3_2 _07654_ (.A(_02075_),
    .B(_02109_),
    .C(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__buf_1 _07655_ (.A(_02112_),
    .X(_00012_));
 sky130_fd_sc_hd__o21ai_2 _07656_ (.A1(\core.mem_do_rdata ),
    .A2(\core.mem_do_wdata ),
    .B1(_02048_),
    .Y(_02113_));
 sky130_fd_sc_hd__a22o_2 _07657_ (.A1(_02079_),
    .A2(_02018_),
    .B1(_02029_),
    .B2(\core.cpu_state[3] ),
    .X(_02114_));
 sky130_fd_sc_hd__inv_2 _07658_ (.A(_02100_),
    .Y(_02115_));
 sky130_fd_sc_hd__buf_1 _07659_ (.A(\core.cpu_state[4] ),
    .X(_02116_));
 sky130_fd_sc_hd__inv_2 _07660_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .Y(_02117_));
 sky130_fd_sc_hd__a22o_2 _07661_ (.A1(_02117_),
    .A2(\core.cpu_state[3] ),
    .B1(\core.cpu_state[1] ),
    .B2(_02108_),
    .X(_02118_));
 sky130_fd_sc_hd__a221o_2 _07662_ (.A1(\core.cpu_state[2] ),
    .A2(_02057_),
    .B1(_02115_),
    .B2(_02116_),
    .C1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__nor2_2 _07663_ (.A(\core.cpu_state[6] ),
    .B(\core.cpu_state[5] ),
    .Y(_02120_));
 sky130_fd_sc_hd__buf_1 _07664_ (.A(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__nor2_2 _07665_ (.A(_02121_),
    .B(_02086_),
    .Y(_00509_));
 sky130_fd_sc_hd__a211o_2 _07666_ (.A1(_02113_),
    .A2(_02114_),
    .B1(_02119_),
    .C1(_00509_),
    .X(_02122_));
 sky130_fd_sc_hd__a21o_2 _07667_ (.A1(_02075_),
    .A2(_02122_),
    .B1(_02055_),
    .X(_00011_));
 sky130_fd_sc_hd__buf_1 _07668_ (.A(_02069_),
    .X(_02123_));
 sky130_fd_sc_hd__o211a_2 _07669_ (.A1(\core.instr_lh ),
    .A2(\core.instr_lhu ),
    .B1(_02051_),
    .C1(_02052_),
    .X(_02124_));
 sky130_fd_sc_hd__a221o_2 _07670_ (.A1(_02123_),
    .A2(_02047_),
    .B1(_02050_),
    .B2(\core.instr_sh ),
    .C1(_02124_),
    .X(_00019_));
 sky130_fd_sc_hd__inv_2 _07671_ (.A(\core.cpu_state[4] ),
    .Y(_02125_));
 sky130_fd_sc_hd__buf_1 _07672_ (.A(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__buf_1 _07673_ (.A(_00004_),
    .X(_02127_));
 sky130_fd_sc_hd__inv_2 _07674_ (.A(_00003_),
    .Y(_02128_));
 sky130_fd_sc_hd__buf_1 _07675_ (.A(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__inv_2 _07676_ (.A(_00002_),
    .Y(_02130_));
 sky130_fd_sc_hd__buf_1 _07677_ (.A(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__buf_1 _07678_ (.A(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__buf_1 _07679_ (.A(_00000_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_1 _07680_ (.A(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_1 _07681_ (.A(_00001_),
    .X(_02135_));
 sky130_fd_sc_hd__mux4_2 _07682_ (.A0(\core.cpuregs[4][2] ),
    .A1(\core.cpuregs[5][2] ),
    .A2(\core.cpuregs[6][2] ),
    .A3(\core.cpuregs[7][2] ),
    .S0(_02134_),
    .S1(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__or2_2 _07683_ (.A(_02132_),
    .B(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__buf_1 _07684_ (.A(_00002_),
    .X(_02138_));
 sky130_fd_sc_hd__buf_1 _07685_ (.A(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_1 _07686_ (.A(_02133_),
    .X(_02140_));
 sky130_fd_sc_hd__mux4_2 _07687_ (.A0(\core.cpuregs[0][2] ),
    .A1(\core.cpuregs[1][2] ),
    .A2(\core.cpuregs[2][2] ),
    .A3(\core.cpuregs[3][2] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_02141_));
 sky130_fd_sc_hd__or2_2 _07688_ (.A(_02139_),
    .B(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__buf_1 _07689_ (.A(_02138_),
    .X(_02143_));
 sky130_fd_sc_hd__buf_1 _07690_ (.A(_00001_),
    .X(_02144_));
 sky130_fd_sc_hd__mux4_2 _07691_ (.A0(\core.cpuregs[8][2] ),
    .A1(\core.cpuregs[9][2] ),
    .A2(\core.cpuregs[10][2] ),
    .A3(\core.cpuregs[11][2] ),
    .S0(_02140_),
    .S1(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__or2_2 _07692_ (.A(_02143_),
    .B(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__buf_1 _07693_ (.A(_02131_),
    .X(_02147_));
 sky130_fd_sc_hd__buf_1 _07694_ (.A(_00000_),
    .X(_02148_));
 sky130_fd_sc_hd__buf_1 _07695_ (.A(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__mux4_2 _07696_ (.A0(\core.cpuregs[12][2] ),
    .A1(\core.cpuregs[13][2] ),
    .A2(\core.cpuregs[14][2] ),
    .A3(\core.cpuregs[15][2] ),
    .S0(_02149_),
    .S1(_02144_),
    .X(_02150_));
 sky130_fd_sc_hd__buf_1 _07697_ (.A(_00003_),
    .X(_02151_));
 sky130_fd_sc_hd__buf_1 _07698_ (.A(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__o21a_2 _07699_ (.A1(_02147_),
    .A2(_02150_),
    .B1(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__a32o_2 _07700_ (.A1(_02129_),
    .A2(_02137_),
    .A3(_02142_),
    .B1(_02146_),
    .B2(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__buf_1 _07701_ (.A(_00000_),
    .X(_02155_));
 sky130_fd_sc_hd__buf_1 _07702_ (.A(_00001_),
    .X(_02156_));
 sky130_fd_sc_hd__mux4_2 _07703_ (.A0(\core.cpuregs[24][2] ),
    .A1(\core.cpuregs[25][2] ),
    .A2(\core.cpuregs[26][2] ),
    .A3(\core.cpuregs[27][2] ),
    .S0(_02155_),
    .S1(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_1 _07704_ (.A(_00001_),
    .X(_02158_));
 sky130_fd_sc_hd__buf_1 _07705_ (.A(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_2 _07706_ (.A0(\core.cpuregs[30][2] ),
    .A1(\core.cpuregs[31][2] ),
    .S(_02148_),
    .X(_02160_));
 sky130_fd_sc_hd__inv_2 _07707_ (.A(_00001_),
    .Y(_02161_));
 sky130_fd_sc_hd__mux2_2 _07708_ (.A0(\core.cpuregs[28][2] ),
    .A1(\core.cpuregs[29][2] ),
    .S(_02133_),
    .X(_02162_));
 sky130_fd_sc_hd__a21o_2 _07709_ (.A1(_02161_),
    .A2(_02162_),
    .B1(_02131_),
    .X(_02163_));
 sky130_fd_sc_hd__a21o_2 _07710_ (.A1(_02159_),
    .A2(_02160_),
    .B1(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__o211a_2 _07711_ (.A1(_02139_),
    .A2(_02157_),
    .B1(_02164_),
    .C1(_02151_),
    .X(_02165_));
 sky130_fd_sc_hd__mux4_2 _07712_ (.A0(\core.cpuregs[20][2] ),
    .A1(\core.cpuregs[21][2] ),
    .A2(\core.cpuregs[22][2] ),
    .A3(\core.cpuregs[23][2] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_02166_));
 sky130_fd_sc_hd__buf_1 _07713_ (.A(_02161_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_2 _07714_ (.A0(\core.cpuregs[16][2] ),
    .A1(\core.cpuregs[17][2] ),
    .S(_02155_),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_2 _07715_ (.A0(\core.cpuregs[18][2] ),
    .A1(\core.cpuregs[19][2] ),
    .S(_02133_),
    .X(_02169_));
 sky130_fd_sc_hd__a21o_2 _07716_ (.A1(_02158_),
    .A2(_02169_),
    .B1(_02138_),
    .X(_02170_));
 sky130_fd_sc_hd__a21o_2 _07717_ (.A1(_02167_),
    .A2(_02168_),
    .B1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__o211a_2 _07718_ (.A1(_02132_),
    .A2(_02166_),
    .B1(_02171_),
    .C1(_02128_),
    .X(_02172_));
 sky130_fd_sc_hd__or3b_2 _07719_ (.A(_02165_),
    .B(_02172_),
    .C_N(_00004_),
    .X(_02173_));
 sky130_fd_sc_hd__or3_2 _07720_ (.A(\core.decoded_imm_j[3] ),
    .B(\core.decoded_imm_j[4] ),
    .C(\core.decoded_imm_j[11] ),
    .X(_02174_));
 sky130_fd_sc_hd__or3_2 _07721_ (.A(\core.decoded_imm_j[1] ),
    .B(\core.decoded_imm_j[2] ),
    .C(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__o211a_2 _07722_ (.A1(_02127_),
    .A2(_02154_),
    .B1(_02173_),
    .C1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__mux2_2 _07723_ (.A0(_02176_),
    .A1(\core.decoded_imm_j[2] ),
    .S(\core.is_slli_srli_srai ),
    .X(_02177_));
 sky130_fd_sc_hd__nor3_2 _07724_ (.A(\core.reg_sh[4] ),
    .B(\core.reg_sh[3] ),
    .C(\core.reg_sh[2] ),
    .Y(_02178_));
 sky130_fd_sc_hd__buf_1 _07725_ (.A(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__o21ai_2 _07726_ (.A1(\core.reg_sh[0] ),
    .A2(\core.reg_sh[1] ),
    .B1(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_2 _07727_ (.A(_02126_),
    .B(\core.reg_sh[2] ),
    .Y(_02181_));
 sky130_fd_sc_hd__a22o_2 _07728_ (.A1(_02126_),
    .A2(_02177_),
    .B1(_02180_),
    .B2(_02181_),
    .X(_00034_));
 sky130_fd_sc_hd__or3b_2 _07729_ (.A(\core.reg_sh[3] ),
    .B(\core.reg_sh[2] ),
    .C_N(\core.reg_sh[4] ),
    .X(_02182_));
 sky130_fd_sc_hd__a21bo_2 _07730_ (.A1(\core.reg_sh[3] ),
    .A2(\core.reg_sh[2] ),
    .B1_N(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__mux4_2 _07731_ (.A0(\core.cpuregs[4][3] ),
    .A1(\core.cpuregs[5][3] ),
    .A2(\core.cpuregs[6][3] ),
    .A3(\core.cpuregs[7][3] ),
    .S0(_02134_),
    .S1(_02135_),
    .X(_02184_));
 sky130_fd_sc_hd__or2_2 _07732_ (.A(_02132_),
    .B(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__mux4_2 _07733_ (.A0(\core.cpuregs[0][3] ),
    .A1(\core.cpuregs[1][3] ),
    .A2(\core.cpuregs[2][3] ),
    .A3(\core.cpuregs[3][3] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_02186_));
 sky130_fd_sc_hd__or2_2 _07734_ (.A(_02139_),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__mux4_2 _07735_ (.A0(\core.cpuregs[8][3] ),
    .A1(\core.cpuregs[9][3] ),
    .A2(\core.cpuregs[10][3] ),
    .A3(\core.cpuregs[11][3] ),
    .S0(_02140_),
    .S1(_02144_),
    .X(_02188_));
 sky130_fd_sc_hd__or2_2 _07736_ (.A(_02143_),
    .B(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__mux4_2 _07737_ (.A0(\core.cpuregs[12][3] ),
    .A1(\core.cpuregs[13][3] ),
    .A2(\core.cpuregs[14][3] ),
    .A3(\core.cpuregs[15][3] ),
    .S0(_02149_),
    .S1(_02144_),
    .X(_02190_));
 sky130_fd_sc_hd__o21a_2 _07738_ (.A1(_02147_),
    .A2(_02190_),
    .B1(_02151_),
    .X(_02191_));
 sky130_fd_sc_hd__a32o_2 _07739_ (.A1(_02128_),
    .A2(_02185_),
    .A3(_02187_),
    .B1(_02189_),
    .B2(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__mux4_2 _07740_ (.A0(\core.cpuregs[24][3] ),
    .A1(\core.cpuregs[25][3] ),
    .A2(\core.cpuregs[26][3] ),
    .A3(\core.cpuregs[27][3] ),
    .S0(_02155_),
    .S1(_02156_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_2 _07741_ (.A0(\core.cpuregs[30][3] ),
    .A1(\core.cpuregs[31][3] ),
    .S(_02148_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_2 _07742_ (.A0(\core.cpuregs[28][3] ),
    .A1(\core.cpuregs[29][3] ),
    .S(_02133_),
    .X(_02195_));
 sky130_fd_sc_hd__a21o_2 _07743_ (.A1(_02161_),
    .A2(_02195_),
    .B1(_02131_),
    .X(_02196_));
 sky130_fd_sc_hd__a21o_2 _07744_ (.A1(_02159_),
    .A2(_02194_),
    .B1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__o211a_2 _07745_ (.A1(_02139_),
    .A2(_02193_),
    .B1(_02197_),
    .C1(_02151_),
    .X(_02198_));
 sky130_fd_sc_hd__mux4_2 _07746_ (.A0(\core.cpuregs[20][3] ),
    .A1(\core.cpuregs[21][3] ),
    .A2(\core.cpuregs[22][3] ),
    .A3(\core.cpuregs[23][3] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_2 _07747_ (.A0(\core.cpuregs[16][3] ),
    .A1(\core.cpuregs[17][3] ),
    .S(_02148_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_2 _07748_ (.A0(\core.cpuregs[18][3] ),
    .A1(\core.cpuregs[19][3] ),
    .S(_02133_),
    .X(_02201_));
 sky130_fd_sc_hd__a21o_2 _07749_ (.A1(_02158_),
    .A2(_02201_),
    .B1(_02138_),
    .X(_02202_));
 sky130_fd_sc_hd__a21o_2 _07750_ (.A1(_02161_),
    .A2(_02200_),
    .B1(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__o211a_2 _07751_ (.A1(_02132_),
    .A2(_02199_),
    .B1(_02203_),
    .C1(_02128_),
    .X(_02204_));
 sky130_fd_sc_hd__or3b_2 _07752_ (.A(_02198_),
    .B(_02204_),
    .C_N(_00004_),
    .X(_02205_));
 sky130_fd_sc_hd__o211a_2 _07753_ (.A1(_02127_),
    .A2(_02192_),
    .B1(_02205_),
    .C1(_02175_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_2 _07754_ (.A0(_02206_),
    .A1(\core.decoded_imm_j[3] ),
    .S(\core.is_slli_srli_srai ),
    .X(_02207_));
 sky130_fd_sc_hd__buf_1 _07755_ (.A(_02116_),
    .X(_02208_));
 sky130_fd_sc_hd__o22a_2 _07756_ (.A1(_02101_),
    .A2(_02183_),
    .B1(_02207_),
    .B2(_02208_),
    .X(_00035_));
 sky130_fd_sc_hd__o21a_2 _07757_ (.A1(\core.reg_sh[3] ),
    .A2(\core.reg_sh[2] ),
    .B1(\core.reg_sh[4] ),
    .X(_02209_));
 sky130_fd_sc_hd__mux4_2 _07758_ (.A0(\core.cpuregs[4][4] ),
    .A1(\core.cpuregs[5][4] ),
    .A2(\core.cpuregs[6][4] ),
    .A3(\core.cpuregs[7][4] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_02210_));
 sky130_fd_sc_hd__or2_2 _07759_ (.A(_02132_),
    .B(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__mux4_2 _07760_ (.A0(\core.cpuregs[0][4] ),
    .A1(\core.cpuregs[1][4] ),
    .A2(\core.cpuregs[2][4] ),
    .A3(\core.cpuregs[3][4] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_02212_));
 sky130_fd_sc_hd__or2_2 _07761_ (.A(_02139_),
    .B(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__mux4_2 _07762_ (.A0(\core.cpuregs[8][4] ),
    .A1(\core.cpuregs[9][4] ),
    .A2(\core.cpuregs[10][4] ),
    .A3(\core.cpuregs[11][4] ),
    .S0(_02140_),
    .S1(_02144_),
    .X(_02214_));
 sky130_fd_sc_hd__or2_2 _07763_ (.A(_02143_),
    .B(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__mux4_2 _07764_ (.A0(\core.cpuregs[12][4] ),
    .A1(\core.cpuregs[13][4] ),
    .A2(\core.cpuregs[14][4] ),
    .A3(\core.cpuregs[15][4] ),
    .S0(_02149_),
    .S1(_02144_),
    .X(_02216_));
 sky130_fd_sc_hd__o21a_2 _07765_ (.A1(_02132_),
    .A2(_02216_),
    .B1(_02151_),
    .X(_02217_));
 sky130_fd_sc_hd__a32o_2 _07766_ (.A1(_02128_),
    .A2(_02211_),
    .A3(_02213_),
    .B1(_02215_),
    .B2(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__mux4_2 _07767_ (.A0(\core.cpuregs[24][4] ),
    .A1(\core.cpuregs[25][4] ),
    .A2(\core.cpuregs[26][4] ),
    .A3(\core.cpuregs[27][4] ),
    .S0(_02155_),
    .S1(_02156_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_2 _07768_ (.A0(\core.cpuregs[30][4] ),
    .A1(\core.cpuregs[31][4] ),
    .S(_02148_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_2 _07769_ (.A0(\core.cpuregs[28][4] ),
    .A1(\core.cpuregs[29][4] ),
    .S(_02133_),
    .X(_02221_));
 sky130_fd_sc_hd__a21o_2 _07770_ (.A1(_02161_),
    .A2(_02221_),
    .B1(_02131_),
    .X(_02222_));
 sky130_fd_sc_hd__a21o_2 _07771_ (.A1(_02144_),
    .A2(_02220_),
    .B1(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__o211a_2 _07772_ (.A1(_02139_),
    .A2(_02219_),
    .B1(_02223_),
    .C1(_02151_),
    .X(_02224_));
 sky130_fd_sc_hd__mux4_2 _07773_ (.A0(\core.cpuregs[20][4] ),
    .A1(\core.cpuregs[21][4] ),
    .A2(\core.cpuregs[22][4] ),
    .A3(\core.cpuregs[23][4] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_2 _07774_ (.A0(\core.cpuregs[16][4] ),
    .A1(\core.cpuregs[17][4] ),
    .S(_02148_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_2 _07775_ (.A0(\core.cpuregs[18][4] ),
    .A1(\core.cpuregs[19][4] ),
    .S(_02133_),
    .X(_02227_));
 sky130_fd_sc_hd__a21o_2 _07776_ (.A1(_02158_),
    .A2(_02227_),
    .B1(_02138_),
    .X(_02228_));
 sky130_fd_sc_hd__a21o_2 _07777_ (.A1(_02161_),
    .A2(_02226_),
    .B1(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__o211a_2 _07778_ (.A1(_02131_),
    .A2(_02225_),
    .B1(_02229_),
    .C1(_02128_),
    .X(_02230_));
 sky130_fd_sc_hd__or3b_2 _07779_ (.A(_02224_),
    .B(_02230_),
    .C_N(_00004_),
    .X(_02231_));
 sky130_fd_sc_hd__o211a_2 _07780_ (.A1(_00004_),
    .A2(_02218_),
    .B1(_02231_),
    .C1(_02175_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_2 _07781_ (.A0(_02232_),
    .A1(\core.decoded_imm_j[4] ),
    .S(\core.is_slli_srli_srai ),
    .X(_02233_));
 sky130_fd_sc_hd__o22a_2 _07782_ (.A1(_02101_),
    .A2(_02209_),
    .B1(_02233_),
    .B2(_02208_),
    .X(_00036_));
 sky130_fd_sc_hd__inv_2 _07783_ (.A(\core.cpu_state[3] ),
    .Y(_02234_));
 sky130_fd_sc_hd__buf_1 _07784_ (.A(_02042_),
    .X(_02235_));
 sky130_fd_sc_hd__buf_1 _07785_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .X(_02236_));
 sky130_fd_sc_hd__buf_1 _07786_ (.A(\core.pcpi_rs1[31] ),
    .X(_02237_));
 sky130_fd_sc_hd__nand2_2 _07787_ (.A(\core.pcpi_rs2[31] ),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__or2_2 _07788_ (.A(\core.pcpi_rs2[31] ),
    .B(\core.pcpi_rs1[31] ),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_2 _07789_ (.A(_02238_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__and2_2 _07790_ (.A(\core.pcpi_rs2[30] ),
    .B(\core.pcpi_rs1[30] ),
    .X(_02241_));
 sky130_fd_sc_hd__buf_1 _07791_ (.A(\core.pcpi_rs1[30] ),
    .X(_02242_));
 sky130_fd_sc_hd__nor2_2 _07792_ (.A(\core.pcpi_rs2[30] ),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__or2_2 _07793_ (.A(_02241_),
    .B(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__and2_2 _07794_ (.A(\core.pcpi_rs2[28] ),
    .B(\core.pcpi_rs1[28] ),
    .X(_02245_));
 sky130_fd_sc_hd__buf_1 _07795_ (.A(\core.pcpi_rs1[28] ),
    .X(_02246_));
 sky130_fd_sc_hd__nor2_2 _07796_ (.A(\core.pcpi_rs2[28] ),
    .B(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__or2_2 _07797_ (.A(_02245_),
    .B(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__and2_2 _07798_ (.A(\core.pcpi_rs2[29] ),
    .B(\core.pcpi_rs1[29] ),
    .X(_02249_));
 sky130_fd_sc_hd__nor2_2 _07799_ (.A(\core.pcpi_rs2[29] ),
    .B(\core.pcpi_rs1[29] ),
    .Y(_02250_));
 sky130_fd_sc_hd__or2_2 _07800_ (.A(_02249_),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__nand4_2 _07801_ (.A(_02240_),
    .B(_02244_),
    .C(_02248_),
    .D(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_2 _07802_ (.A(\core.pcpi_rs2[25] ),
    .B(\core.pcpi_rs1[25] ),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_2 _07803_ (.A(\core.pcpi_rs2[25] ),
    .B(\core.pcpi_rs1[25] ),
    .Y(_02254_));
 sky130_fd_sc_hd__nand2b_2 _07804_ (.A_N(_02253_),
    .B(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__buf_1 _07805_ (.A(\core.pcpi_rs1[24] ),
    .X(_02256_));
 sky130_fd_sc_hd__nor2_2 _07806_ (.A(\core.pcpi_rs2[24] ),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_2 _07807_ (.A(\core.pcpi_rs2[24] ),
    .B(\core.pcpi_rs1[24] ),
    .Y(_02258_));
 sky130_fd_sc_hd__nand2b_2 _07808_ (.A_N(_02257_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__nand2_2 _07809_ (.A(_02255_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__and2_2 _07810_ (.A(\core.pcpi_rs2[27] ),
    .B(\core.pcpi_rs1[27] ),
    .X(_02261_));
 sky130_fd_sc_hd__nor2_2 _07811_ (.A(\core.pcpi_rs2[27] ),
    .B(\core.pcpi_rs1[27] ),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_2 _07812_ (.A(_02261_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__and2_2 _07813_ (.A(\core.pcpi_rs2[26] ),
    .B(\core.pcpi_rs1[26] ),
    .X(_02264_));
 sky130_fd_sc_hd__nor2_2 _07814_ (.A(\core.pcpi_rs2[26] ),
    .B(\core.pcpi_rs1[26] ),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_2 _07815_ (.A(_02264_),
    .B(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__or3_2 _07816_ (.A(_02260_),
    .B(_02263_),
    .C(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__nor2_2 _07817_ (.A(_02252_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__and2_2 _07818_ (.A(\core.pcpi_rs2[23] ),
    .B(\core.pcpi_rs1[23] ),
    .X(_02269_));
 sky130_fd_sc_hd__buf_1 _07819_ (.A(\core.pcpi_rs1[23] ),
    .X(_02270_));
 sky130_fd_sc_hd__nor2_2 _07820_ (.A(\core.pcpi_rs2[23] ),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__or2_2 _07821_ (.A(_02269_),
    .B(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__and2_2 _07822_ (.A(\core.pcpi_rs2[22] ),
    .B(\core.pcpi_rs1[22] ),
    .X(_02273_));
 sky130_fd_sc_hd__nor2_2 _07823_ (.A(\core.pcpi_rs2[22] ),
    .B(\core.pcpi_rs1[22] ),
    .Y(_02274_));
 sky130_fd_sc_hd__or2_2 _07824_ (.A(_02273_),
    .B(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__or2_2 _07825_ (.A(\core.pcpi_rs2[20] ),
    .B(\core.pcpi_rs1[20] ),
    .X(_02276_));
 sky130_fd_sc_hd__buf_1 _07826_ (.A(\core.pcpi_rs1[20] ),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_2 _07827_ (.A(\core.pcpi_rs2[20] ),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_2 _07828_ (.A(_02276_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_2 _07829_ (.A(\core.pcpi_rs2[21] ),
    .B(\core.pcpi_rs1[21] ),
    .Y(_02280_));
 sky130_fd_sc_hd__buf_1 _07830_ (.A(\core.pcpi_rs1[21] ),
    .X(_02281_));
 sky130_fd_sc_hd__nand2_2 _07831_ (.A(\core.pcpi_rs2[21] ),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand2b_2 _07832_ (.A_N(_02280_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand4_2 _07833_ (.A(_02272_),
    .B(_02275_),
    .C(_02279_),
    .D(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__inv_2 _07834_ (.A(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__xor2_2 _07835_ (.A(\core.pcpi_rs2[19] ),
    .B(\core.pcpi_rs1[19] ),
    .X(_02286_));
 sky130_fd_sc_hd__nor2_2 _07836_ (.A(\core.pcpi_rs2[18] ),
    .B(\core.pcpi_rs1[18] ),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_2 _07837_ (.A(\core.pcpi_rs2[18] ),
    .B(\core.pcpi_rs1[18] ),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2b_2 _07838_ (.A_N(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__inv_2 _07839_ (.A(\core.pcpi_rs2[16] ),
    .Y(_02290_));
 sky130_fd_sc_hd__buf_1 _07840_ (.A(\core.pcpi_rs1[16] ),
    .X(_02291_));
 sky130_fd_sc_hd__or2_2 _07841_ (.A(\core.pcpi_rs2[17] ),
    .B(\core.pcpi_rs1[17] ),
    .X(_02292_));
 sky130_fd_sc_hd__buf_1 _07842_ (.A(\core.pcpi_rs1[17] ),
    .X(_02293_));
 sky130_fd_sc_hd__nand2_2 _07843_ (.A(\core.pcpi_rs2[17] ),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_2 _07844_ (.A(_02292_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__and2b_2 _07845_ (.A_N(\core.pcpi_rs2[17] ),
    .B(_02293_),
    .X(_02296_));
 sky130_fd_sc_hd__a31o_2 _07846_ (.A1(_02290_),
    .A2(_02291_),
    .A3(_02295_),
    .B1(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__buf_1 _07847_ (.A(\core.pcpi_rs1[18] ),
    .X(_02298_));
 sky130_fd_sc_hd__and2b_2 _07848_ (.A_N(\core.pcpi_rs2[18] ),
    .B(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__a21oi_2 _07849_ (.A1(_02289_),
    .A2(_02297_),
    .B1(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__inv_2 _07850_ (.A(\core.pcpi_rs2[15] ),
    .Y(_02301_));
 sky130_fd_sc_hd__inv_2 _07851_ (.A(\core.pcpi_rs1[15] ),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_2 _07852_ (.A(_02301_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_2 _07853_ (.A(\core.pcpi_rs2[15] ),
    .B(\core.pcpi_rs1[15] ),
    .Y(_02304_));
 sky130_fd_sc_hd__or2_2 _07854_ (.A(_02303_),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__buf_1 _07855_ (.A(\core.pcpi_rs1[14] ),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_2 _07856_ (.A(\core.pcpi_rs2[14] ),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor2_2 _07857_ (.A(\core.pcpi_rs2[14] ),
    .B(\core.pcpi_rs1[14] ),
    .Y(_02308_));
 sky130_fd_sc_hd__inv_2 _07858_ (.A(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__nand2_2 _07859_ (.A(_02307_),
    .B(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_2 _07860_ (.A(\core.pcpi_rs2[13] ),
    .B(\core.pcpi_rs1[13] ),
    .Y(_02311_));
 sky130_fd_sc_hd__buf_1 _07861_ (.A(\core.pcpi_rs1[13] ),
    .X(_02312_));
 sky130_fd_sc_hd__nand2_2 _07862_ (.A(\core.pcpi_rs2[13] ),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2b_2 _07863_ (.A_N(_02311_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__buf_1 _07864_ (.A(\core.pcpi_rs1[12] ),
    .X(_02315_));
 sky130_fd_sc_hd__nor2_2 _07865_ (.A(\core.pcpi_rs2[12] ),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__nand2_2 _07866_ (.A(\core.pcpi_rs2[12] ),
    .B(\core.pcpi_rs1[12] ),
    .Y(_02317_));
 sky130_fd_sc_hd__nand2b_2 _07867_ (.A_N(_02316_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__and2_2 _07868_ (.A(\core.pcpi_rs2[11] ),
    .B(\core.pcpi_rs1[11] ),
    .X(_02319_));
 sky130_fd_sc_hd__nor2_2 _07869_ (.A(\core.pcpi_rs2[11] ),
    .B(\core.pcpi_rs1[11] ),
    .Y(_02320_));
 sky130_fd_sc_hd__or2_2 _07870_ (.A(_02319_),
    .B(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__or2_2 _07871_ (.A(\core.pcpi_rs2[10] ),
    .B(\core.pcpi_rs1[10] ),
    .X(_02322_));
 sky130_fd_sc_hd__buf_1 _07872_ (.A(\core.pcpi_rs1[10] ),
    .X(_02323_));
 sky130_fd_sc_hd__nand2_2 _07873_ (.A(\core.pcpi_rs2[10] ),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_2 _07874_ (.A(_02322_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__inv_2 _07875_ (.A(\core.pcpi_rs2[8] ),
    .Y(_02326_));
 sky130_fd_sc_hd__buf_1 _07876_ (.A(\core.pcpi_rs1[8] ),
    .X(_02327_));
 sky130_fd_sc_hd__nor2_2 _07877_ (.A(\core.pcpi_rs2[9] ),
    .B(\core.pcpi_rs1[9] ),
    .Y(_02328_));
 sky130_fd_sc_hd__nand2_2 _07878_ (.A(\core.pcpi_rs2[9] ),
    .B(\core.pcpi_rs1[9] ),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2b_2 _07879_ (.A_N(_02328_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__buf_1 _07880_ (.A(\core.pcpi_rs1[9] ),
    .X(_02331_));
 sky130_fd_sc_hd__and2b_2 _07881_ (.A_N(\core.pcpi_rs2[9] ),
    .B(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__a31o_2 _07882_ (.A1(_02326_),
    .A2(_02327_),
    .A3(_02330_),
    .B1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__and2b_2 _07883_ (.A_N(\core.pcpi_rs2[10] ),
    .B(_02323_),
    .X(_02334_));
 sky130_fd_sc_hd__a21o_2 _07884_ (.A1(_02325_),
    .A2(_02333_),
    .B1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__buf_1 _07885_ (.A(\core.pcpi_rs1[11] ),
    .X(_02336_));
 sky130_fd_sc_hd__and2b_2 _07886_ (.A_N(\core.pcpi_rs2[11] ),
    .B(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__a21o_2 _07887_ (.A1(_02321_),
    .A2(_02335_),
    .B1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__inv_2 _07888_ (.A(\core.pcpi_rs2[12] ),
    .Y(_02339_));
 sky130_fd_sc_hd__and2b_2 _07889_ (.A_N(\core.pcpi_rs2[13] ),
    .B(_02312_),
    .X(_02340_));
 sky130_fd_sc_hd__a31o_2 _07890_ (.A1(_02339_),
    .A2(_02315_),
    .A3(_02314_),
    .B1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__a31o_2 _07891_ (.A1(_02314_),
    .A2(_02318_),
    .A3(_02338_),
    .B1(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__and2b_2 _07892_ (.A_N(\core.pcpi_rs2[14] ),
    .B(_02306_),
    .X(_02343_));
 sky130_fd_sc_hd__a21o_2 _07893_ (.A1(_02310_),
    .A2(_02342_),
    .B1(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__buf_1 _07894_ (.A(\core.pcpi_rs1[15] ),
    .X(_02345_));
 sky130_fd_sc_hd__or2_2 _07895_ (.A(\core.pcpi_rs2[8] ),
    .B(\core.pcpi_rs1[8] ),
    .X(_02346_));
 sky130_fd_sc_hd__nand2_2 _07896_ (.A(\core.pcpi_rs2[8] ),
    .B(\core.pcpi_rs1[8] ),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_2 _07897_ (.A(_02346_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__and4_2 _07898_ (.A(_02321_),
    .B(_02325_),
    .C(_02330_),
    .D(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__and3_2 _07899_ (.A(_02310_),
    .B(_02314_),
    .C(_02318_),
    .X(_02350_));
 sky130_fd_sc_hd__and3_2 _07900_ (.A(_02305_),
    .B(_02349_),
    .C(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__nor2_2 _07901_ (.A(\core.mem_la_wdata[5] ),
    .B(\core.pcpi_rs1[5] ),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_2 _07902_ (.A(\core.mem_la_wdata[5] ),
    .B(\core.pcpi_rs1[5] ),
    .Y(_02353_));
 sky130_fd_sc_hd__or2b_2 _07903_ (.A(_02352_),
    .B_N(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_1 _07904_ (.A(\core.pcpi_rs1[4] ),
    .X(_02355_));
 sky130_fd_sc_hd__and2_2 _07905_ (.A(\core.mem_la_wdata[4] ),
    .B(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__nor2_2 _07906_ (.A(\core.mem_la_wdata[4] ),
    .B(\core.pcpi_rs1[4] ),
    .Y(_02357_));
 sky130_fd_sc_hd__or2_2 _07907_ (.A(_02356_),
    .B(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__nand2_2 _07908_ (.A(\core.mem_la_wdata[3] ),
    .B(\core.pcpi_rs1[3] ),
    .Y(_02359_));
 sky130_fd_sc_hd__or2_2 _07909_ (.A(\core.mem_la_wdata[3] ),
    .B(\core.pcpi_rs1[3] ),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_2 _07910_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_2 _07911_ (.A(\core.mem_la_wdata[2] ),
    .B(\core.pcpi_rs1[2] ),
    .Y(_02362_));
 sky130_fd_sc_hd__or2_2 _07912_ (.A(\core.mem_la_wdata[2] ),
    .B(\core.pcpi_rs1[2] ),
    .X(_02363_));
 sky130_fd_sc_hd__nand2_2 _07913_ (.A(_02362_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__inv_2 _07914_ (.A(_02071_),
    .Y(_02365_));
 sky130_fd_sc_hd__buf_1 _07915_ (.A(\core.mem_la_wdata[1] ),
    .X(_02366_));
 sky130_fd_sc_hd__inv_2 _07916_ (.A(\core.pcpi_rs1[0] ),
    .Y(_02367_));
 sky130_fd_sc_hd__buf_1 _07917_ (.A(\core.mem_la_wdata[0] ),
    .X(_02368_));
 sky130_fd_sc_hd__xor2_2 _07918_ (.A(\core.pcpi_rs1[1] ),
    .B(_02366_),
    .X(_02369_));
 sky130_fd_sc_hd__a21oi_2 _07919_ (.A1(_02367_),
    .A2(_02368_),
    .B1(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__o21bai_2 _07920_ (.A1(_02365_),
    .A2(_02366_),
    .B1_N(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__buf_1 _07921_ (.A(\core.pcpi_rs1[2] ),
    .X(_02372_));
 sky130_fd_sc_hd__and2b_2 _07922_ (.A_N(\core.mem_la_wdata[2] ),
    .B(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__a21o_2 _07923_ (.A1(_02364_),
    .A2(_02371_),
    .B1(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__buf_1 _07924_ (.A(\core.pcpi_rs1[3] ),
    .X(_02375_));
 sky130_fd_sc_hd__and2b_2 _07925_ (.A_N(\core.mem_la_wdata[3] ),
    .B(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__a21o_2 _07926_ (.A1(_02361_),
    .A2(_02374_),
    .B1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__and3_2 _07927_ (.A(_02354_),
    .B(_02358_),
    .C(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__and2_2 _07928_ (.A(\core.mem_la_wdata[7] ),
    .B(\core.pcpi_rs1[7] ),
    .X(_02379_));
 sky130_fd_sc_hd__buf_1 _07929_ (.A(\core.pcpi_rs1[7] ),
    .X(_02380_));
 sky130_fd_sc_hd__nor2_2 _07930_ (.A(\core.mem_la_wdata[7] ),
    .B(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__or2_2 _07931_ (.A(_02379_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__buf_1 _07932_ (.A(\core.pcpi_rs1[6] ),
    .X(_02383_));
 sky130_fd_sc_hd__nand2_2 _07933_ (.A(\core.mem_la_wdata[6] ),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__or2_2 _07934_ (.A(\core.mem_la_wdata[6] ),
    .B(\core.pcpi_rs1[6] ),
    .X(_02385_));
 sky130_fd_sc_hd__nand2_2 _07935_ (.A(_02384_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__inv_2 _07936_ (.A(\core.mem_la_wdata[4] ),
    .Y(_02387_));
 sky130_fd_sc_hd__buf_1 _07937_ (.A(\core.pcpi_rs1[5] ),
    .X(_02388_));
 sky130_fd_sc_hd__and2b_2 _07938_ (.A_N(\core.mem_la_wdata[5] ),
    .B(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__a31o_2 _07939_ (.A1(_02387_),
    .A2(_02355_),
    .A3(_02354_),
    .B1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__and2b_2 _07940_ (.A_N(\core.mem_la_wdata[6] ),
    .B(_02383_),
    .X(_02391_));
 sky130_fd_sc_hd__a21o_2 _07941_ (.A1(_02386_),
    .A2(_02390_),
    .B1(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__and2b_2 _07942_ (.A_N(\core.mem_la_wdata[7] ),
    .B(_02380_),
    .X(_02393_));
 sky130_fd_sc_hd__a21o_2 _07943_ (.A1(_02382_),
    .A2(_02392_),
    .B1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__a31o_2 _07944_ (.A1(_02378_),
    .A2(_02382_),
    .A3(_02386_),
    .B1(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__a22o_2 _07945_ (.A1(_02301_),
    .A2(_02345_),
    .B1(_02351_),
    .B2(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__a21oi_2 _07946_ (.A1(_02305_),
    .A2(_02344_),
    .B1(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__nor2_2 _07947_ (.A(\core.pcpi_rs2[16] ),
    .B(_02291_),
    .Y(_02398_));
 sky130_fd_sc_hd__and2_2 _07948_ (.A(\core.pcpi_rs2[16] ),
    .B(\core.pcpi_rs1[16] ),
    .X(_02399_));
 sky130_fd_sc_hd__nor2_2 _07949_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_2 _07950_ (.A(_02289_),
    .B(_02295_),
    .Y(_02401_));
 sky130_fd_sc_hd__or3_2 _07951_ (.A(_02286_),
    .B(_02400_),
    .C(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__or2b_2 _07952_ (.A(\core.pcpi_rs2[19] ),
    .B_N(\core.pcpi_rs1[19] ),
    .X(_02403_));
 sky130_fd_sc_hd__o221ai_2 _07953_ (.A1(_02286_),
    .A2(_02300_),
    .B1(_02397_),
    .B2(_02402_),
    .C1(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__inv_2 _07954_ (.A(\core.pcpi_rs2[20] ),
    .Y(_02405_));
 sky130_fd_sc_hd__and2b_2 _07955_ (.A_N(\core.pcpi_rs2[21] ),
    .B(_02281_),
    .X(_02406_));
 sky130_fd_sc_hd__a31o_2 _07956_ (.A1(_02405_),
    .A2(_02277_),
    .A3(_02283_),
    .B1(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__buf_1 _07957_ (.A(\core.pcpi_rs1[22] ),
    .X(_02408_));
 sky130_fd_sc_hd__and2b_2 _07958_ (.A_N(\core.pcpi_rs2[22] ),
    .B(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__a21o_2 _07959_ (.A1(_02275_),
    .A2(_02407_),
    .B1(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__and2b_2 _07960_ (.A_N(\core.pcpi_rs2[23] ),
    .B(_02270_),
    .X(_02411_));
 sky130_fd_sc_hd__a221o_2 _07961_ (.A1(_02285_),
    .A2(_02404_),
    .B1(_02410_),
    .B2(_02272_),
    .C1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__and2b_2 _07962_ (.A_N(\core.pcpi_rs2[28] ),
    .B(_02246_),
    .X(_02413_));
 sky130_fd_sc_hd__buf_1 _07963_ (.A(\core.pcpi_rs1[29] ),
    .X(_02414_));
 sky130_fd_sc_hd__and2b_2 _07964_ (.A_N(\core.pcpi_rs2[29] ),
    .B(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__a21o_2 _07965_ (.A1(_02251_),
    .A2(_02413_),
    .B1(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__and2b_2 _07966_ (.A_N(\core.pcpi_rs2[30] ),
    .B(_02242_),
    .X(_02417_));
 sky130_fd_sc_hd__a21o_2 _07967_ (.A1(_02244_),
    .A2(_02416_),
    .B1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__and2b_2 _07968_ (.A_N(\core.pcpi_rs2[24] ),
    .B(_02256_),
    .X(_02419_));
 sky130_fd_sc_hd__and2b_2 _07969_ (.A_N(\core.pcpi_rs2[25] ),
    .B(\core.pcpi_rs1[25] ),
    .X(_02420_));
 sky130_fd_sc_hd__a21oi_2 _07970_ (.A1(_02255_),
    .A2(_02419_),
    .B1(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__buf_1 _07971_ (.A(\core.pcpi_rs1[26] ),
    .X(_02422_));
 sky130_fd_sc_hd__or2b_2 _07972_ (.A(\core.pcpi_rs2[26] ),
    .B_N(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__o21a_2 _07973_ (.A1(_02266_),
    .A2(_02421_),
    .B1(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__or2b_2 _07974_ (.A(\core.pcpi_rs2[27] ),
    .B_N(\core.pcpi_rs1[27] ),
    .X(_02425_));
 sky130_fd_sc_hd__o21a_2 _07975_ (.A1(_02263_),
    .A2(_02424_),
    .B1(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__nor2_2 _07976_ (.A(_02252_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__a221o_2 _07977_ (.A1(_02268_),
    .A2(_02412_),
    .B1(_02418_),
    .B2(_02240_),
    .C1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__and2b_2 _07978_ (.A_N(\core.pcpi_rs2[31] ),
    .B(_02237_),
    .X(_02429_));
 sky130_fd_sc_hd__nor2_2 _07979_ (.A(_02428_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__o21a_2 _07980_ (.A1(_02428_),
    .A2(_02429_),
    .B1(\core.instr_bgeu ),
    .X(_02431_));
 sky130_fd_sc_hd__nor4_2 _07981_ (.A(\core.instr_bne ),
    .B(\core.is_slti_blt_slt ),
    .C(\core.is_sltiu_bltu_sltu ),
    .D(_02058_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_2 _07982_ (.A(_02361_),
    .B(_02364_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_2 _07983_ (.A(_02070_),
    .B(_02368_),
    .Y(_02434_));
 sky130_fd_sc_hd__or2_2 _07984_ (.A(\core.pcpi_rs1[0] ),
    .B(_02368_),
    .X(_02435_));
 sky130_fd_sc_hd__and2_2 _07985_ (.A(_02434_),
    .B(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__and4_2 _07986_ (.A(_02354_),
    .B(_02358_),
    .C(_02382_),
    .D(_02386_),
    .X(_02437_));
 sky130_fd_sc_hd__or4b_2 _07987_ (.A(_02369_),
    .B(_02433_),
    .C(_02436_),
    .D_N(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_2 _07988_ (.A(_02268_),
    .B(_02351_),
    .Y(_02439_));
 sky130_fd_sc_hd__or4_2 _07989_ (.A(_02284_),
    .B(_02402_),
    .C(_02438_),
    .D(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_2 _07990_ (.A0(_02432_),
    .A1(\core.instr_bne ),
    .S(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__inv_2 _07991_ (.A(_02428_),
    .Y(_02442_));
 sky130_fd_sc_hd__a21o_2 _07992_ (.A1(_02240_),
    .A2(_02442_),
    .B1(_02429_),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_2 _07993_ (.A0(\core.instr_bge ),
    .A1(\core.is_slti_blt_slt ),
    .S(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__a2111o_2 _07994_ (.A1(\core.is_sltiu_bltu_sltu ),
    .A2(_02430_),
    .B1(_02431_),
    .C1(_02441_),
    .D1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_2 _07995_ (.A(_02236_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__and3_2 _07996_ (.A(\core.mem_do_rinst ),
    .B(resetn),
    .C(_02029_),
    .X(_02447_));
 sky130_fd_sc_hd__buf_1 _07997_ (.A(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__buf_1 _07998_ (.A(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__o32a_2 _07999_ (.A1(_02234_),
    .A2(_02235_),
    .A3(_02446_),
    .B1(_02449_),
    .B2(_00509_),
    .X(_00030_));
 sky130_fd_sc_hd__buf_1 _08000_ (.A(\core.cpu_state[3] ),
    .X(_02450_));
 sky130_fd_sc_hd__buf_1 _08001_ (.A(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__and3_2 _08002_ (.A(_02234_),
    .B(_02126_),
    .C(_02036_),
    .X(_02452_));
 sky130_fd_sc_hd__buf_1 _08003_ (.A(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__buf_1 _08004_ (.A(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__buf_1 _08005_ (.A(\core.instr_rdinstrh ),
    .X(_02455_));
 sky130_fd_sc_hd__buf_1 _08006_ (.A(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__nor3_2 _08007_ (.A(\core.instr_rdinstr ),
    .B(\core.instr_rdinstrh ),
    .C(\core.instr_rdcycleh ),
    .Y(_02457_));
 sky130_fd_sc_hd__buf_1 _08008_ (.A(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__buf_1 _08009_ (.A(\core.instr_rdinstr ),
    .X(_02459_));
 sky130_fd_sc_hd__buf_1 _08010_ (.A(\core.instr_rdcycleh ),
    .X(_02460_));
 sky130_fd_sc_hd__a22o_2 _08011_ (.A1(\core.count_instr[0] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[32] ),
    .X(_02461_));
 sky130_fd_sc_hd__a221o_2 _08012_ (.A1(\core.count_instr[32] ),
    .A2(_02456_),
    .B1(_02458_),
    .B2(\core.count_cycle[0] ),
    .C1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__buf_1 _08013_ (.A(_02116_),
    .X(_02463_));
 sky130_fd_sc_hd__nor2_2 _08014_ (.A(\core.mem_wordsize[1] ),
    .B(\core.mem_wordsize[2] ),
    .Y(_02464_));
 sky130_fd_sc_hd__a21o_2 _08015_ (.A1(\core.mem_wordsize[2] ),
    .A2(_02365_),
    .B1(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2b_2 _08016_ (.A_N(_02465_),
    .B(_02072_),
    .Y(_02466_));
 sky130_fd_sc_hd__and2_2 _08017_ (.A(\core.mem_wordsize[1] ),
    .B(_02070_),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_2 _08018_ (.A0(mem_rdata[8]),
    .A1(mem_rdata[24]),
    .S(_02071_),
    .X(_02468_));
 sky130_fd_sc_hd__o21a_2 _08019_ (.A1(\core.mem_wordsize[2] ),
    .A2(_02367_),
    .B1(_02071_),
    .X(_02469_));
 sky130_fd_sc_hd__a22o_2 _08020_ (.A1(_02467_),
    .A2(_02468_),
    .B1(_02469_),
    .B2(mem_rdata[16]),
    .X(_02470_));
 sky130_fd_sc_hd__or2_2 _08021_ (.A(_02023_),
    .B(\core.mem_wordsize[2] ),
    .X(_02471_));
 sky130_fd_sc_hd__buf_1 _08022_ (.A(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__a22o_2 _08023_ (.A1(mem_rdata[0]),
    .A2(_02466_),
    .B1(_02470_),
    .B2(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__a22o_2 _08024_ (.A1(_02463_),
    .A2(_02070_),
    .B1(_02473_),
    .B2(_02087_),
    .X(_02474_));
 sky130_fd_sc_hd__a221o_2 _08025_ (.A1(_02451_),
    .A2(\core.decoded_imm[0] ),
    .B1(_02454_),
    .B2(_02462_),
    .C1(_02474_),
    .X(_01543_));
 sky130_fd_sc_hd__buf_1 _08026_ (.A(_02071_),
    .X(_02475_));
 sky130_fd_sc_hd__buf_1 _08027_ (.A(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_2 _08028_ (.A0(mem_rdata[9]),
    .A1(mem_rdata[25]),
    .S(_02475_),
    .X(_02477_));
 sky130_fd_sc_hd__a22o_2 _08029_ (.A1(mem_rdata[17]),
    .A2(_02469_),
    .B1(_02477_),
    .B2(_02467_),
    .X(_02478_));
 sky130_fd_sc_hd__a22o_2 _08030_ (.A1(mem_rdata[1]),
    .A2(_02466_),
    .B1(_02478_),
    .B2(_02472_),
    .X(_02479_));
 sky130_fd_sc_hd__buf_1 _08031_ (.A(_02045_),
    .X(_02480_));
 sky130_fd_sc_hd__nand2_2 _08032_ (.A(\core.reg_pc[1] ),
    .B(\core.decoded_imm[1] ),
    .Y(_02481_));
 sky130_fd_sc_hd__or2_2 _08033_ (.A(\core.reg_pc[1] ),
    .B(\core.decoded_imm[1] ),
    .X(_02482_));
 sky130_fd_sc_hd__and3_2 _08034_ (.A(\core.cpu_state[3] ),
    .B(_02481_),
    .C(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__a221o_2 _08035_ (.A1(_02463_),
    .A2(_02476_),
    .B1(_02479_),
    .B2(_02480_),
    .C1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__buf_1 _08036_ (.A(_02458_),
    .X(_02485_));
 sky130_fd_sc_hd__buf_1 _08037_ (.A(\core.instr_rdinstrh ),
    .X(_02486_));
 sky130_fd_sc_hd__or3_2 _08038_ (.A(\core.cpu_state[3] ),
    .B(\core.cpu_state[4] ),
    .C(\core.cpu_state[6] ),
    .X(_02487_));
 sky130_fd_sc_hd__buf_1 _08039_ (.A(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__buf_1 _08040_ (.A(\core.instr_rdcycleh ),
    .X(_02489_));
 sky130_fd_sc_hd__a22o_2 _08041_ (.A1(\core.count_instr[1] ),
    .A2(_02459_),
    .B1(_02489_),
    .B2(\core.count_cycle[33] ),
    .X(_02490_));
 sky130_fd_sc_hd__a211o_2 _08042_ (.A1(\core.count_instr[33] ),
    .A2(_02486_),
    .B1(_02488_),
    .C1(_02490_),
    .X(_02491_));
 sky130_fd_sc_hd__a21o_2 _08043_ (.A1(\core.count_cycle[1] ),
    .A2(_02485_),
    .B1(_02491_),
    .X(_02492_));
 sky130_fd_sc_hd__o21a_2 _08044_ (.A1(_02454_),
    .A2(_02484_),
    .B1(_02492_),
    .X(_01554_));
 sky130_fd_sc_hd__buf_1 _08045_ (.A(\core.reg_pc[2] ),
    .X(_02493_));
 sky130_fd_sc_hd__xor2_2 _08046_ (.A(_02493_),
    .B(\core.decoded_imm[2] ),
    .X(_02494_));
 sky130_fd_sc_hd__xnor2_2 _08047_ (.A(_02481_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__a22o_2 _08048_ (.A1(_02116_),
    .A2(_02372_),
    .B1(_02495_),
    .B2(_02450_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_2 _08049_ (.A0(mem_rdata[10]),
    .A1(mem_rdata[26]),
    .S(_02071_),
    .X(_02497_));
 sky130_fd_sc_hd__a22o_2 _08050_ (.A1(mem_rdata[18]),
    .A2(_02469_),
    .B1(_02497_),
    .B2(_02467_),
    .X(_02498_));
 sky130_fd_sc_hd__a22o_2 _08051_ (.A1(mem_rdata[2]),
    .A2(_02466_),
    .B1(_02498_),
    .B2(_02472_),
    .X(_02499_));
 sky130_fd_sc_hd__a22o_2 _08052_ (.A1(\core.count_instr[2] ),
    .A2(\core.instr_rdinstr ),
    .B1(\core.instr_rdcycleh ),
    .B2(\core.count_cycle[34] ),
    .X(_02500_));
 sky130_fd_sc_hd__a221o_2 _08053_ (.A1(\core.count_instr[34] ),
    .A2(_02455_),
    .B1(\core.count_cycle[2] ),
    .B2(_02457_),
    .C1(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__a22o_2 _08054_ (.A1(_02045_),
    .A2(_02499_),
    .B1(_02501_),
    .B2(_02453_),
    .X(_02502_));
 sky130_fd_sc_hd__or2_2 _08055_ (.A(_02496_),
    .B(_02502_),
    .X(_02503_));
 sky130_fd_sc_hd__buf_1 _08056_ (.A(_02503_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_2 _08057_ (.A0(mem_rdata[11]),
    .A1(mem_rdata[27]),
    .S(_02475_),
    .X(_02504_));
 sky130_fd_sc_hd__a22o_2 _08058_ (.A1(mem_rdata[19]),
    .A2(_02469_),
    .B1(_02504_),
    .B2(_02467_),
    .X(_02505_));
 sky130_fd_sc_hd__a22o_2 _08059_ (.A1(mem_rdata[3]),
    .A2(_02466_),
    .B1(_02505_),
    .B2(_02472_),
    .X(_02506_));
 sky130_fd_sc_hd__a22o_2 _08060_ (.A1(\core.reg_pc[1] ),
    .A2(\core.decoded_imm[1] ),
    .B1(\core.decoded_imm[2] ),
    .B2(_02493_),
    .X(_02507_));
 sky130_fd_sc_hd__o21ai_2 _08061_ (.A1(_02493_),
    .A2(\core.decoded_imm[2] ),
    .B1(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__nand2_2 _08062_ (.A(\core.reg_pc[3] ),
    .B(\core.decoded_imm[3] ),
    .Y(_02509_));
 sky130_fd_sc_hd__inv_2 _08063_ (.A(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_2 _08064_ (.A(\core.reg_pc[3] ),
    .B(\core.decoded_imm[3] ),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_2 _08065_ (.A(_02510_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__xnor2_2 _08066_ (.A(_02508_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__buf_1 _08067_ (.A(_02453_),
    .X(_02514_));
 sky130_fd_sc_hd__buf_1 _08068_ (.A(\core.instr_rdinstr ),
    .X(_02515_));
 sky130_fd_sc_hd__a22o_2 _08069_ (.A1(\core.count_instr[3] ),
    .A2(_02515_),
    .B1(_02489_),
    .B2(\core.count_cycle[35] ),
    .X(_02516_));
 sky130_fd_sc_hd__a221o_2 _08070_ (.A1(\core.count_instr[35] ),
    .A2(_02455_),
    .B1(\core.count_cycle[3] ),
    .B2(_02458_),
    .C1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__a22o_2 _08071_ (.A1(_02463_),
    .A2(_02375_),
    .B1(_02514_),
    .B2(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__a221o_2 _08072_ (.A1(_02480_),
    .A2(_02506_),
    .B1(_02513_),
    .B2(_02451_),
    .C1(_02518_),
    .X(_01568_));
 sky130_fd_sc_hd__a21o_2 _08073_ (.A1(_02508_),
    .A2(_02509_),
    .B1(_02511_),
    .X(_02519_));
 sky130_fd_sc_hd__or2_2 _08074_ (.A(\core.reg_pc[4] ),
    .B(\core.decoded_imm[4] ),
    .X(_02520_));
 sky130_fd_sc_hd__nand2_2 _08075_ (.A(\core.reg_pc[4] ),
    .B(\core.decoded_imm[4] ),
    .Y(_02521_));
 sky130_fd_sc_hd__nand2_2 _08076_ (.A(_02520_),
    .B(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__buf_1 _08077_ (.A(\core.cpu_state[3] ),
    .X(_02523_));
 sky130_fd_sc_hd__o21ai_2 _08078_ (.A1(_02519_),
    .A2(_02522_),
    .B1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__a21oi_2 _08079_ (.A1(_02519_),
    .A2(_02522_),
    .B1(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__mux2_2 _08080_ (.A0(mem_rdata[12]),
    .A1(mem_rdata[28]),
    .S(_02475_),
    .X(_02526_));
 sky130_fd_sc_hd__a22o_2 _08081_ (.A1(mem_rdata[20]),
    .A2(_02469_),
    .B1(_02526_),
    .B2(_02467_),
    .X(_02527_));
 sky130_fd_sc_hd__a22o_2 _08082_ (.A1(mem_rdata[4]),
    .A2(_02466_),
    .B1(_02527_),
    .B2(_02472_),
    .X(_02528_));
 sky130_fd_sc_hd__a221o_2 _08083_ (.A1(_02463_),
    .A2(_02355_),
    .B1(_02528_),
    .B2(_02087_),
    .C1(_02514_),
    .X(_02529_));
 sky130_fd_sc_hd__buf_1 _08084_ (.A(_02458_),
    .X(_02530_));
 sky130_fd_sc_hd__buf_1 _08085_ (.A(_02488_),
    .X(_02531_));
 sky130_fd_sc_hd__buf_1 _08086_ (.A(_02489_),
    .X(_02532_));
 sky130_fd_sc_hd__a22o_2 _08087_ (.A1(\core.count_instr[4] ),
    .A2(_02515_),
    .B1(_02455_),
    .B2(\core.count_instr[36] ),
    .X(_02533_));
 sky130_fd_sc_hd__a21o_2 _08088_ (.A1(_02532_),
    .A2(\core.count_cycle[36] ),
    .B1(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__a211o_2 _08089_ (.A1(\core.count_cycle[4] ),
    .A2(_02530_),
    .B1(_02531_),
    .C1(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__o21a_2 _08090_ (.A1(_02525_),
    .A2(_02529_),
    .B1(_02535_),
    .X(_01569_));
 sky130_fd_sc_hd__a22o_2 _08091_ (.A1(\core.count_instr[5] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[37] ),
    .X(_02536_));
 sky130_fd_sc_hd__a211o_2 _08092_ (.A1(\core.count_instr[37] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__a21oi_2 _08093_ (.A1(\core.count_cycle[5] ),
    .A2(_02485_),
    .B1(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__or2_2 _08094_ (.A(\core.reg_pc[5] ),
    .B(\core.decoded_imm[5] ),
    .X(_02539_));
 sky130_fd_sc_hd__nand2_2 _08095_ (.A(\core.reg_pc[5] ),
    .B(\core.decoded_imm[5] ),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_2 _08096_ (.A(_02539_),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__o21a_2 _08097_ (.A1(_02519_),
    .A2(_02522_),
    .B1(_02521_),
    .X(_02542_));
 sky130_fd_sc_hd__nand2_2 _08098_ (.A(_02541_),
    .B(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21a_2 _08099_ (.A1(_02541_),
    .A2(_02542_),
    .B1(_02450_),
    .X(_02544_));
 sky130_fd_sc_hd__buf_1 _08100_ (.A(\core.cpu_state[4] ),
    .X(_02545_));
 sky130_fd_sc_hd__buf_1 _08101_ (.A(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_2 _08102_ (.A0(mem_rdata[13]),
    .A1(mem_rdata[29]),
    .S(_02071_),
    .X(_02547_));
 sky130_fd_sc_hd__a22o_2 _08103_ (.A1(mem_rdata[21]),
    .A2(_02469_),
    .B1(_02547_),
    .B2(_02467_),
    .X(_02548_));
 sky130_fd_sc_hd__a22o_2 _08104_ (.A1(mem_rdata[5]),
    .A2(_02466_),
    .B1(_02548_),
    .B2(_02472_),
    .X(_02549_));
 sky130_fd_sc_hd__a221o_2 _08105_ (.A1(_02546_),
    .A2(_02388_),
    .B1(_02549_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02550_));
 sky130_fd_sc_hd__a21oi_2 _08106_ (.A1(_02543_),
    .A2(_02544_),
    .B1(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2_2 _08107_ (.A(_02538_),
    .B(_02551_),
    .Y(_01570_));
 sky130_fd_sc_hd__a22o_2 _08108_ (.A1(\core.count_instr[6] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[38] ),
    .X(_02552_));
 sky130_fd_sc_hd__a211o_2 _08109_ (.A1(\core.count_instr[38] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__a21oi_2 _08110_ (.A1(\core.count_cycle[6] ),
    .A2(_02485_),
    .B1(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand3_2 _08111_ (.A(\core.reg_pc[4] ),
    .B(\core.decoded_imm[4] ),
    .C(_02539_),
    .Y(_02555_));
 sky130_fd_sc_hd__or3_2 _08112_ (.A(_02519_),
    .B(_02522_),
    .C(_02541_),
    .X(_02556_));
 sky130_fd_sc_hd__and3_2 _08113_ (.A(_02540_),
    .B(_02555_),
    .C(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__or2_2 _08114_ (.A(\core.reg_pc[6] ),
    .B(\core.decoded_imm[6] ),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_2 _08115_ (.A(\core.reg_pc[6] ),
    .B(\core.decoded_imm[6] ),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_2 _08116_ (.A(_02558_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__xor2_2 _08117_ (.A(_02557_),
    .B(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_2 _08118_ (.A0(mem_rdata[14]),
    .A1(mem_rdata[30]),
    .S(_02071_),
    .X(_02562_));
 sky130_fd_sc_hd__a22o_2 _08119_ (.A1(mem_rdata[22]),
    .A2(_02469_),
    .B1(_02562_),
    .B2(_02467_),
    .X(_02563_));
 sky130_fd_sc_hd__a22o_2 _08120_ (.A1(mem_rdata[6]),
    .A2(_02466_),
    .B1(_02563_),
    .B2(_02472_),
    .X(_02564_));
 sky130_fd_sc_hd__a221o_2 _08121_ (.A1(_02546_),
    .A2(_02383_),
    .B1(_02564_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02565_));
 sky130_fd_sc_hd__a21oi_2 _08122_ (.A1(_02451_),
    .A2(_02561_),
    .B1(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_2 _08123_ (.A(_02554_),
    .B(_02566_),
    .Y(_01571_));
 sky130_fd_sc_hd__a22o_2 _08124_ (.A1(\core.count_instr[7] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[39] ),
    .X(_02567_));
 sky130_fd_sc_hd__a211o_2 _08125_ (.A1(\core.count_instr[39] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__a21oi_2 _08126_ (.A1(\core.count_cycle[7] ),
    .A2(_02485_),
    .B1(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__or2_2 _08127_ (.A(\core.reg_pc[7] ),
    .B(\core.decoded_imm[7] ),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_2 _08128_ (.A(\core.reg_pc[7] ),
    .B(\core.decoded_imm[7] ),
    .Y(_02571_));
 sky130_fd_sc_hd__nand2_2 _08129_ (.A(_02570_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__o21ai_2 _08130_ (.A1(_02557_),
    .A2(_02560_),
    .B1(_02559_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_2 _08131_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__mux2_2 _08132_ (.A0(mem_rdata[15]),
    .A1(mem_rdata[31]),
    .S(_02071_),
    .X(_02575_));
 sky130_fd_sc_hd__a22o_2 _08133_ (.A1(mem_rdata[23]),
    .A2(_02469_),
    .B1(_02575_),
    .B2(_02467_),
    .X(_02576_));
 sky130_fd_sc_hd__a22o_2 _08134_ (.A1(mem_rdata[7]),
    .A2(_02466_),
    .B1(_02576_),
    .B2(_02472_),
    .X(_02577_));
 sky130_fd_sc_hd__a221o_2 _08135_ (.A1(_02546_),
    .A2(_02380_),
    .B1(_02577_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02578_));
 sky130_fd_sc_hd__a21oi_2 _08136_ (.A1(_02523_),
    .A2(_02574_),
    .B1(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__nor2_2 _08137_ (.A(_02569_),
    .B(_02579_),
    .Y(_01572_));
 sky130_fd_sc_hd__and3_2 _08138_ (.A(\core.reg_pc[6] ),
    .B(\core.decoded_imm[6] ),
    .C(_02570_),
    .X(_02580_));
 sky130_fd_sc_hd__a21oi_2 _08139_ (.A1(\core.reg_pc[7] ),
    .A2(\core.decoded_imm[7] ),
    .B1(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__a311o_2 _08140_ (.A1(_02540_),
    .A2(_02555_),
    .A3(_02556_),
    .B1(_02560_),
    .C1(_02572_),
    .X(_02582_));
 sky130_fd_sc_hd__and2_2 _08141_ (.A(_02581_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__or2_2 _08142_ (.A(\core.reg_pc[8] ),
    .B(\core.decoded_imm[8] ),
    .X(_02584_));
 sky130_fd_sc_hd__nand2_2 _08143_ (.A(\core.reg_pc[8] ),
    .B(\core.decoded_imm[8] ),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_2 _08144_ (.A(_02584_),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__xor2_2 _08145_ (.A(_02583_),
    .B(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__or2b_2 _08146_ (.A(\core.latched_is_lh ),
    .B_N(\core.latched_is_lb ),
    .X(_02588_));
 sky130_fd_sc_hd__a32o_2 _08147_ (.A1(_02123_),
    .A2(_02476_),
    .A3(mem_rdata[24]),
    .B1(_02465_),
    .B2(mem_rdata[8]),
    .X(_02589_));
 sky130_fd_sc_hd__and2_2 _08148_ (.A(\core.latched_is_lb ),
    .B(_02577_),
    .X(_02590_));
 sky130_fd_sc_hd__a21o_2 _08149_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__a22o_2 _08150_ (.A1(\core.count_instr[8] ),
    .A2(_02515_),
    .B1(_02489_),
    .B2(\core.count_cycle[40] ),
    .X(_02592_));
 sky130_fd_sc_hd__a221o_2 _08151_ (.A1(\core.count_instr[40] ),
    .A2(_02455_),
    .B1(\core.count_cycle[8] ),
    .B2(_02458_),
    .C1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__a22o_2 _08152_ (.A1(_02463_),
    .A2(_02327_),
    .B1(_02514_),
    .B2(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__a221o_2 _08153_ (.A1(_02451_),
    .A2(_02587_),
    .B1(_02591_),
    .B2(_02480_),
    .C1(_02594_),
    .X(_01573_));
 sky130_fd_sc_hd__a22o_2 _08154_ (.A1(\core.count_instr[9] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[41] ),
    .X(_02595_));
 sky130_fd_sc_hd__a211o_2 _08155_ (.A1(\core.count_instr[41] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__a21oi_2 _08156_ (.A1(\core.count_cycle[9] ),
    .A2(_02485_),
    .B1(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_2 _08157_ (.A(\core.reg_pc[9] ),
    .B(\core.decoded_imm[9] ),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_2 _08158_ (.A(\core.reg_pc[9] ),
    .B(\core.decoded_imm[9] ),
    .Y(_02599_));
 sky130_fd_sc_hd__nand2_2 _08159_ (.A(_02598_),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__o21a_2 _08160_ (.A1(_02583_),
    .A2(_02586_),
    .B1(_02585_),
    .X(_02601_));
 sky130_fd_sc_hd__nand2_2 _08161_ (.A(_02600_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__o21a_2 _08162_ (.A1(_02600_),
    .A2(_02601_),
    .B1(_02450_),
    .X(_02603_));
 sky130_fd_sc_hd__a32o_2 _08163_ (.A1(_02069_),
    .A2(_02475_),
    .A3(mem_rdata[25]),
    .B1(_02465_),
    .B2(mem_rdata[9]),
    .X(_02604_));
 sky130_fd_sc_hd__a21o_2 _08164_ (.A1(_02588_),
    .A2(_02604_),
    .B1(_02590_),
    .X(_02605_));
 sky130_fd_sc_hd__a221o_2 _08165_ (.A1(_02546_),
    .A2(_02331_),
    .B1(_02605_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02606_));
 sky130_fd_sc_hd__a21oi_2 _08166_ (.A1(_02602_),
    .A2(_02603_),
    .B1(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nor2_2 _08167_ (.A(_02597_),
    .B(_02607_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand3_2 _08168_ (.A(\core.reg_pc[8] ),
    .B(\core.decoded_imm[8] ),
    .C(_02598_),
    .Y(_02608_));
 sky130_fd_sc_hd__a211o_2 _08169_ (.A1(_02581_),
    .A2(_02582_),
    .B1(_02586_),
    .C1(_02600_),
    .X(_02609_));
 sky130_fd_sc_hd__nand3_2 _08170_ (.A(_02599_),
    .B(_02608_),
    .C(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hd__or2_2 _08171_ (.A(\core.reg_pc[10] ),
    .B(\core.decoded_imm[10] ),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_2 _08172_ (.A(\core.reg_pc[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_02612_));
 sky130_fd_sc_hd__nand2_2 _08173_ (.A(_02611_),
    .B(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__xnor2_2 _08174_ (.A(_02610_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a32o_2 _08175_ (.A1(_02123_),
    .A2(_02476_),
    .A3(mem_rdata[26]),
    .B1(_02465_),
    .B2(mem_rdata[10]),
    .X(_02615_));
 sky130_fd_sc_hd__a21o_2 _08176_ (.A1(_02588_),
    .A2(_02615_),
    .B1(_02590_),
    .X(_02616_));
 sky130_fd_sc_hd__a22o_2 _08177_ (.A1(\core.count_instr[10] ),
    .A2(\core.instr_rdinstr ),
    .B1(\core.instr_rdcycleh ),
    .B2(\core.count_cycle[42] ),
    .X(_02617_));
 sky130_fd_sc_hd__a221o_2 _08178_ (.A1(\core.count_instr[42] ),
    .A2(_02455_),
    .B1(\core.count_cycle[10] ),
    .B2(_02457_),
    .C1(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a22o_2 _08179_ (.A1(_02463_),
    .A2(_02323_),
    .B1(_02514_),
    .B2(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__a221o_2 _08180_ (.A1(_02451_),
    .A2(_02614_),
    .B1(_02616_),
    .B2(_02480_),
    .C1(_02619_),
    .X(_01544_));
 sky130_fd_sc_hd__a22o_2 _08181_ (.A1(\core.count_instr[11] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[43] ),
    .X(_02620_));
 sky130_fd_sc_hd__a211o_2 _08182_ (.A1(\core.count_instr[43] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_2 _08183_ (.A1(\core.count_cycle[11] ),
    .A2(_02485_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__or2_2 _08184_ (.A(\core.reg_pc[11] ),
    .B(\core.decoded_imm[11] ),
    .X(_02623_));
 sky130_fd_sc_hd__nand2_2 _08185_ (.A(\core.reg_pc[11] ),
    .B(\core.decoded_imm[11] ),
    .Y(_02624_));
 sky130_fd_sc_hd__nand2_2 _08186_ (.A(_02623_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__a21bo_2 _08187_ (.A1(_02610_),
    .A2(_02611_),
    .B1_N(_02612_),
    .X(_02626_));
 sky130_fd_sc_hd__xnor2_2 _08188_ (.A(_02625_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__a32o_2 _08189_ (.A1(_02069_),
    .A2(_02475_),
    .A3(mem_rdata[27]),
    .B1(_02465_),
    .B2(mem_rdata[11]),
    .X(_02628_));
 sky130_fd_sc_hd__a21o_2 _08190_ (.A1(_02588_),
    .A2(_02628_),
    .B1(_02590_),
    .X(_02629_));
 sky130_fd_sc_hd__a221o_2 _08191_ (.A1(_02546_),
    .A2(_02336_),
    .B1(_02629_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02630_));
 sky130_fd_sc_hd__a21oi_2 _08192_ (.A1(_02523_),
    .A2(_02627_),
    .B1(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__nor2_2 _08193_ (.A(_02622_),
    .B(_02631_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand3_2 _08194_ (.A(\core.reg_pc[10] ),
    .B(\core.decoded_imm[10] ),
    .C(_02623_),
    .Y(_02632_));
 sky130_fd_sc_hd__a311o_2 _08195_ (.A1(_02599_),
    .A2(_02608_),
    .A3(_02609_),
    .B1(_02613_),
    .C1(_02625_),
    .X(_02633_));
 sky130_fd_sc_hd__and3_2 _08196_ (.A(_02624_),
    .B(_02632_),
    .C(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__or2_2 _08197_ (.A(\core.reg_pc[12] ),
    .B(\core.decoded_imm[12] ),
    .X(_02635_));
 sky130_fd_sc_hd__nand2_2 _08198_ (.A(\core.reg_pc[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_02636_));
 sky130_fd_sc_hd__nand2_2 _08199_ (.A(_02635_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__xor2_2 _08200_ (.A(_02634_),
    .B(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__a32o_2 _08201_ (.A1(_02123_),
    .A2(_02476_),
    .A3(mem_rdata[28]),
    .B1(_02465_),
    .B2(mem_rdata[12]),
    .X(_02639_));
 sky130_fd_sc_hd__a21o_2 _08202_ (.A1(_02588_),
    .A2(_02639_),
    .B1(_02590_),
    .X(_02640_));
 sky130_fd_sc_hd__a22o_2 _08203_ (.A1(\core.count_instr[12] ),
    .A2(\core.instr_rdinstr ),
    .B1(\core.instr_rdcycleh ),
    .B2(\core.count_cycle[44] ),
    .X(_02641_));
 sky130_fd_sc_hd__a221o_2 _08204_ (.A1(\core.count_instr[44] ),
    .A2(_02455_),
    .B1(\core.count_cycle[12] ),
    .B2(_02457_),
    .C1(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__a22o_2 _08205_ (.A1(_02463_),
    .A2(_02315_),
    .B1(_02514_),
    .B2(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__a221o_2 _08206_ (.A1(_02451_),
    .A2(_02638_),
    .B1(_02640_),
    .B2(_02480_),
    .C1(_02643_),
    .X(_01546_));
 sky130_fd_sc_hd__a22o_2 _08207_ (.A1(\core.count_instr[13] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[45] ),
    .X(_02644_));
 sky130_fd_sc_hd__a211o_2 _08208_ (.A1(\core.count_instr[45] ),
    .A2(_02456_),
    .B1(_02531_),
    .C1(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__a21oi_2 _08209_ (.A1(\core.count_cycle[13] ),
    .A2(_02485_),
    .B1(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__or2_2 _08210_ (.A(\core.reg_pc[13] ),
    .B(\core.decoded_imm[13] ),
    .X(_02647_));
 sky130_fd_sc_hd__nand2_2 _08211_ (.A(\core.reg_pc[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_2 _08212_ (.A(_02647_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__o21ai_2 _08213_ (.A1(_02634_),
    .A2(_02637_),
    .B1(_02636_),
    .Y(_02650_));
 sky130_fd_sc_hd__xnor2_2 _08214_ (.A(_02649_),
    .B(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__a32o_2 _08215_ (.A1(_02069_),
    .A2(_02475_),
    .A3(mem_rdata[29]),
    .B1(_02465_),
    .B2(mem_rdata[13]),
    .X(_02652_));
 sky130_fd_sc_hd__a21o_2 _08216_ (.A1(_02588_),
    .A2(_02652_),
    .B1(_02590_),
    .X(_02653_));
 sky130_fd_sc_hd__a221o_2 _08217_ (.A1(_02546_),
    .A2(_02312_),
    .B1(_02653_),
    .B2(_02087_),
    .C1(_02453_),
    .X(_02654_));
 sky130_fd_sc_hd__a21oi_2 _08218_ (.A1(_02523_),
    .A2(_02651_),
    .B1(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__nor2_2 _08219_ (.A(_02646_),
    .B(_02655_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand3_2 _08220_ (.A(\core.reg_pc[12] ),
    .B(\core.decoded_imm[12] ),
    .C(_02647_),
    .Y(_02656_));
 sky130_fd_sc_hd__a311o_2 _08221_ (.A1(_02624_),
    .A2(_02632_),
    .A3(_02633_),
    .B1(_02637_),
    .C1(_02649_),
    .X(_02657_));
 sky130_fd_sc_hd__and3_2 _08222_ (.A(_02648_),
    .B(_02656_),
    .C(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__or2_2 _08223_ (.A(\core.reg_pc[14] ),
    .B(\core.decoded_imm[14] ),
    .X(_02659_));
 sky130_fd_sc_hd__nand2_2 _08224_ (.A(\core.reg_pc[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2_2 _08225_ (.A(_02659_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__xor2_2 _08226_ (.A(_02658_),
    .B(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__a32o_2 _08227_ (.A1(_02123_),
    .A2(_02476_),
    .A3(mem_rdata[30]),
    .B1(_02465_),
    .B2(mem_rdata[14]),
    .X(_02663_));
 sky130_fd_sc_hd__a21o_2 _08228_ (.A1(_02588_),
    .A2(_02663_),
    .B1(_02590_),
    .X(_02664_));
 sky130_fd_sc_hd__a22o_2 _08229_ (.A1(\core.count_instr[14] ),
    .A2(\core.instr_rdinstr ),
    .B1(\core.instr_rdcycleh ),
    .B2(\core.count_cycle[46] ),
    .X(_02665_));
 sky130_fd_sc_hd__a221o_2 _08230_ (.A1(\core.count_instr[46] ),
    .A2(_02455_),
    .B1(\core.count_cycle[14] ),
    .B2(_02457_),
    .C1(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__a22o_2 _08231_ (.A1(_02463_),
    .A2(_02306_),
    .B1(_02514_),
    .B2(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__a221o_2 _08232_ (.A1(_02451_),
    .A2(_02662_),
    .B1(_02664_),
    .B2(_02480_),
    .C1(_02667_),
    .X(_01548_));
 sky130_fd_sc_hd__a22o_2 _08233_ (.A1(\core.count_instr[15] ),
    .A2(_02459_),
    .B1(_02460_),
    .B2(\core.count_cycle[47] ),
    .X(_02668_));
 sky130_fd_sc_hd__a211o_2 _08234_ (.A1(\core.count_instr[47] ),
    .A2(_02456_),
    .B1(_02488_),
    .C1(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__a21oi_2 _08235_ (.A1(\core.count_cycle[15] ),
    .A2(_02485_),
    .B1(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__xnor2_2 _08236_ (.A(\core.reg_pc[15] ),
    .B(\core.decoded_imm[15] ),
    .Y(_02671_));
 sky130_fd_sc_hd__o21ai_2 _08237_ (.A1(_02658_),
    .A2(_02661_),
    .B1(_02660_),
    .Y(_02672_));
 sky130_fd_sc_hd__xnor2_2 _08238_ (.A(_02671_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__or2_2 _08239_ (.A(\core.latched_is_lh ),
    .B(\core.latched_is_lb ),
    .X(_02674_));
 sky130_fd_sc_hd__buf_1 _08240_ (.A(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__a32o_2 _08241_ (.A1(_02069_),
    .A2(_02071_),
    .A3(mem_rdata[31]),
    .B1(_02465_),
    .B2(mem_rdata[15]),
    .X(_02676_));
 sky130_fd_sc_hd__a21oi_2 _08242_ (.A1(\core.latched_is_lh ),
    .A2(_02676_),
    .B1(_02590_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_2 _08243_ (.A(_02675_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__o211a_2 _08244_ (.A1(_02675_),
    .A2(_02676_),
    .B1(_02678_),
    .C1(_02045_),
    .X(_02679_));
 sky130_fd_sc_hd__a211o_2 _08245_ (.A1(_02463_),
    .A2(_02345_),
    .B1(_02453_),
    .C1(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__a21oi_2 _08246_ (.A1(_02523_),
    .A2(_02673_),
    .B1(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_2 _08247_ (.A(_02670_),
    .B(_02681_),
    .Y(_01549_));
 sky130_fd_sc_hd__buf_1 _08248_ (.A(_02531_),
    .X(_02682_));
 sky130_fd_sc_hd__and2_2 _08249_ (.A(\core.count_instr[48] ),
    .B(_02486_),
    .X(_02683_));
 sky130_fd_sc_hd__buf_1 _08250_ (.A(_02515_),
    .X(_02684_));
 sky130_fd_sc_hd__a22o_2 _08251_ (.A1(\core.count_instr[16] ),
    .A2(_02684_),
    .B1(_02532_),
    .B2(\core.count_cycle[48] ),
    .X(_02685_));
 sky130_fd_sc_hd__a211o_2 _08252_ (.A1(\core.count_cycle[16] ),
    .A2(_02530_),
    .B1(_02683_),
    .C1(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__o211a_2 _08253_ (.A1(\core.reg_pc[15] ),
    .A2(\core.decoded_imm[15] ),
    .B1(\core.decoded_imm[14] ),
    .C1(\core.reg_pc[14] ),
    .X(_02687_));
 sky130_fd_sc_hd__a21oi_2 _08254_ (.A1(\core.reg_pc[15] ),
    .A2(\core.decoded_imm[15] ),
    .B1(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__a311o_2 _08255_ (.A1(_02648_),
    .A2(_02656_),
    .A3(_02657_),
    .B1(_02661_),
    .C1(_02671_),
    .X(_02689_));
 sky130_fd_sc_hd__nand2_2 _08256_ (.A(_02688_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__nor2_2 _08257_ (.A(\core.reg_pc[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_02691_));
 sky130_fd_sc_hd__and2_2 _08258_ (.A(\core.reg_pc[16] ),
    .B(\core.decoded_imm[16] ),
    .X(_02692_));
 sky130_fd_sc_hd__nor2_2 _08259_ (.A(_02691_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__xor2_2 _08260_ (.A(_02690_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__buf_1 _08261_ (.A(_02464_),
    .X(_02695_));
 sky130_fd_sc_hd__a21o_2 _08262_ (.A1(mem_rdata[16]),
    .A2(_02695_),
    .B1(_02675_),
    .X(_02696_));
 sky130_fd_sc_hd__a32o_2 _08263_ (.A1(_02045_),
    .A2(_02678_),
    .A3(_02696_),
    .B1(_02291_),
    .B2(_02116_),
    .X(_02697_));
 sky130_fd_sc_hd__a211o_2 _08264_ (.A1(_02523_),
    .A2(_02694_),
    .B1(_02697_),
    .C1(_02454_),
    .X(_02698_));
 sky130_fd_sc_hd__o21a_2 _08265_ (.A1(_02682_),
    .A2(_02686_),
    .B1(_02698_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_2 _08266_ (.A(\core.reg_pc[17] ),
    .B(\core.decoded_imm[17] ),
    .X(_02699_));
 sky130_fd_sc_hd__nor2_2 _08267_ (.A(\core.reg_pc[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_02700_));
 sky130_fd_sc_hd__nor2_2 _08268_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__a21o_2 _08269_ (.A1(_02690_),
    .A2(_02693_),
    .B1(_02692_),
    .X(_02702_));
 sky130_fd_sc_hd__or2_2 _08270_ (.A(_02701_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__nand2_2 _08271_ (.A(_02701_),
    .B(_02702_),
    .Y(_02704_));
 sky130_fd_sc_hd__a22o_2 _08272_ (.A1(\core.count_instr[17] ),
    .A2(_02515_),
    .B1(\core.instr_rdinstrh ),
    .B2(\core.count_instr[49] ),
    .X(_02705_));
 sky130_fd_sc_hd__a221o_2 _08273_ (.A1(_02460_),
    .A2(\core.count_cycle[49] ),
    .B1(\core.count_cycle[17] ),
    .B2(_02458_),
    .C1(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__nand2_2 _08274_ (.A(_02045_),
    .B(_02678_),
    .Y(_02707_));
 sky130_fd_sc_hd__buf_1 _08275_ (.A(_02464_),
    .X(_02708_));
 sky130_fd_sc_hd__buf_1 _08276_ (.A(_02675_),
    .X(_02709_));
 sky130_fd_sc_hd__a21oi_2 _08277_ (.A1(mem_rdata[17]),
    .A2(_02708_),
    .B1(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_2 _08278_ (.A(_02707_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a221o_2 _08279_ (.A1(_02208_),
    .A2(_02293_),
    .B1(_02514_),
    .B2(_02706_),
    .C1(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__a31o_2 _08280_ (.A1(_02451_),
    .A2(_02703_),
    .A3(_02704_),
    .B1(_02712_),
    .X(_01551_));
 sky130_fd_sc_hd__or2_2 _08281_ (.A(\core.reg_pc[18] ),
    .B(\core.decoded_imm[18] ),
    .X(_02713_));
 sky130_fd_sc_hd__nand2_2 _08282_ (.A(\core.reg_pc[18] ),
    .B(\core.decoded_imm[18] ),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_2 _08283_ (.A(_02713_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__o21bai_2 _08284_ (.A1(_02692_),
    .A2(_02699_),
    .B1_N(_02700_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_2 _08285_ (.A(_02693_),
    .B(_02701_),
    .Y(_02717_));
 sky130_fd_sc_hd__a21o_2 _08286_ (.A1(_02688_),
    .A2(_02689_),
    .B1(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__and3_2 _08287_ (.A(_02715_),
    .B(_02716_),
    .C(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__a21o_2 _08288_ (.A1(_02716_),
    .A2(_02718_),
    .B1(_02715_),
    .X(_02720_));
 sky130_fd_sc_hd__and3b_2 _08289_ (.A_N(_02719_),
    .B(_02720_),
    .C(_02450_),
    .X(_02721_));
 sky130_fd_sc_hd__buf_1 _08290_ (.A(_02464_),
    .X(_02722_));
 sky130_fd_sc_hd__a21o_2 _08291_ (.A1(mem_rdata[18]),
    .A2(_02722_),
    .B1(_02709_),
    .X(_02723_));
 sky130_fd_sc_hd__a32o_2 _08292_ (.A1(_02480_),
    .A2(_02678_),
    .A3(_02723_),
    .B1(_02298_),
    .B2(_02208_),
    .X(_02724_));
 sky130_fd_sc_hd__a22o_2 _08293_ (.A1(\core.count_instr[18] ),
    .A2(_02515_),
    .B1(_02489_),
    .B2(\core.count_cycle[50] ),
    .X(_02725_));
 sky130_fd_sc_hd__a211o_2 _08294_ (.A1(\core.count_instr[50] ),
    .A2(_02486_),
    .B1(_02488_),
    .C1(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__a21o_2 _08295_ (.A1(\core.count_cycle[18] ),
    .A2(_02485_),
    .B1(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__o31a_2 _08296_ (.A1(_02454_),
    .A2(_02721_),
    .A3(_02724_),
    .B1(_02727_),
    .X(_01552_));
 sky130_fd_sc_hd__and2_2 _08297_ (.A(\core.count_instr[51] ),
    .B(_02486_),
    .X(_02728_));
 sky130_fd_sc_hd__a22o_2 _08298_ (.A1(\core.count_instr[19] ),
    .A2(_02684_),
    .B1(_02532_),
    .B2(\core.count_cycle[51] ),
    .X(_02729_));
 sky130_fd_sc_hd__a211o_2 _08299_ (.A1(\core.count_cycle[19] ),
    .A2(_02530_),
    .B1(_02728_),
    .C1(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__or2_2 _08300_ (.A(\core.reg_pc[19] ),
    .B(\core.decoded_imm[19] ),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_2 _08301_ (.A(\core.reg_pc[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_2 _08302_ (.A(_02731_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__a21oi_2 _08303_ (.A1(_02714_),
    .A2(_02720_),
    .B1(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__a31o_2 _08304_ (.A1(_02714_),
    .A2(_02720_),
    .A3(_02733_),
    .B1(_02234_),
    .X(_02735_));
 sky130_fd_sc_hd__buf_1 _08305_ (.A(\core.pcpi_rs1[19] ),
    .X(_02736_));
 sky130_fd_sc_hd__a21oi_2 _08306_ (.A1(mem_rdata[19]),
    .A2(_02695_),
    .B1(_02709_),
    .Y(_02737_));
 sky130_fd_sc_hd__o2bb2a_2 _08307_ (.A1_N(_02546_),
    .A2_N(_02736_),
    .B1(_02707_),
    .B2(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__o211ai_2 _08308_ (.A1(_02734_),
    .A2(_02735_),
    .B1(_02738_),
    .C1(_02682_),
    .Y(_02739_));
 sky130_fd_sc_hd__o21a_2 _08309_ (.A1(_02682_),
    .A2(_02730_),
    .B1(_02739_),
    .X(_01553_));
 sky130_fd_sc_hd__or2_2 _08310_ (.A(\core.reg_pc[20] ),
    .B(\core.decoded_imm[20] ),
    .X(_02740_));
 sky130_fd_sc_hd__nand2_2 _08311_ (.A(\core.reg_pc[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_2 _08312_ (.A(_02740_),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__or2_2 _08313_ (.A(_02715_),
    .B(_02733_),
    .X(_02743_));
 sky130_fd_sc_hd__nor2_2 _08314_ (.A(_02717_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__o21ai_2 _08315_ (.A1(_02716_),
    .A2(_02743_),
    .B1(_02732_),
    .Y(_02745_));
 sky130_fd_sc_hd__a31o_2 _08316_ (.A1(\core.reg_pc[18] ),
    .A2(\core.decoded_imm[18] ),
    .A3(_02731_),
    .B1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a21oi_2 _08317_ (.A1(_02690_),
    .A2(_02744_),
    .B1(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand2_2 _08318_ (.A(_02742_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__or2_2 _08319_ (.A(_02742_),
    .B(_02747_),
    .X(_02749_));
 sky130_fd_sc_hd__and3_2 _08320_ (.A(_02450_),
    .B(_02748_),
    .C(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__a21o_2 _08321_ (.A1(mem_rdata[20]),
    .A2(_02722_),
    .B1(_02709_),
    .X(_02751_));
 sky130_fd_sc_hd__a32o_2 _08322_ (.A1(_02480_),
    .A2(_02678_),
    .A3(_02751_),
    .B1(_02277_),
    .B2(_02208_),
    .X(_02752_));
 sky130_fd_sc_hd__a22o_2 _08323_ (.A1(\core.count_instr[52] ),
    .A2(_02455_),
    .B1(_02489_),
    .B2(\core.count_cycle[52] ),
    .X(_02753_));
 sky130_fd_sc_hd__a211o_2 _08324_ (.A1(\core.count_instr[20] ),
    .A2(_02684_),
    .B1(_02488_),
    .C1(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__a21o_2 _08325_ (.A1(\core.count_cycle[20] ),
    .A2(_02530_),
    .B1(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__o31a_2 _08326_ (.A1(_02454_),
    .A2(_02750_),
    .A3(_02752_),
    .B1(_02755_),
    .X(_01555_));
 sky130_fd_sc_hd__nand2_2 _08327_ (.A(\core.reg_pc[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_02756_));
 sky130_fd_sc_hd__inv_2 _08328_ (.A(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__nor2_2 _08329_ (.A(\core.reg_pc[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_02758_));
 sky130_fd_sc_hd__nor2_2 _08330_ (.A(_02757_),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2_2 _08331_ (.A(_02741_),
    .B(_02749_),
    .Y(_02760_));
 sky130_fd_sc_hd__or2_2 _08332_ (.A(_02759_),
    .B(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__nand2_2 _08333_ (.A(_02759_),
    .B(_02760_),
    .Y(_02762_));
 sky130_fd_sc_hd__a22o_2 _08334_ (.A1(\core.count_instr[21] ),
    .A2(_02515_),
    .B1(\core.instr_rdinstrh ),
    .B2(\core.count_instr[53] ),
    .X(_02763_));
 sky130_fd_sc_hd__a221o_2 _08335_ (.A1(_02460_),
    .A2(\core.count_cycle[53] ),
    .B1(\core.count_cycle[21] ),
    .B2(_02458_),
    .C1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__a21oi_2 _08336_ (.A1(mem_rdata[21]),
    .A2(_02722_),
    .B1(_02709_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_2 _08337_ (.A(_02707_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__a221o_2 _08338_ (.A1(_02208_),
    .A2(_02281_),
    .B1(_02514_),
    .B2(_02764_),
    .C1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__a31o_2 _08339_ (.A1(_02451_),
    .A2(_02761_),
    .A3(_02762_),
    .B1(_02767_),
    .X(_01556_));
 sky130_fd_sc_hd__and2_2 _08340_ (.A(\core.count_instr[54] ),
    .B(_02486_),
    .X(_02768_));
 sky130_fd_sc_hd__a22o_2 _08341_ (.A1(\core.count_instr[22] ),
    .A2(_02684_),
    .B1(_02532_),
    .B2(\core.count_cycle[54] ),
    .X(_02769_));
 sky130_fd_sc_hd__a211o_2 _08342_ (.A1(\core.count_cycle[22] ),
    .A2(_02530_),
    .B1(_02768_),
    .C1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__nor2_2 _08343_ (.A(_02757_),
    .B(_02760_),
    .Y(_02771_));
 sky130_fd_sc_hd__or2_2 _08344_ (.A(\core.reg_pc[22] ),
    .B(\core.decoded_imm[22] ),
    .X(_02772_));
 sky130_fd_sc_hd__nand2_2 _08345_ (.A(\core.reg_pc[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_2 _08346_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o21ai_2 _08347_ (.A1(_02758_),
    .A2(_02771_),
    .B1(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__or3_2 _08348_ (.A(_02758_),
    .B(_02774_),
    .C(_02771_),
    .X(_02776_));
 sky130_fd_sc_hd__a21o_2 _08349_ (.A1(mem_rdata[22]),
    .A2(_02464_),
    .B1(_02675_),
    .X(_02777_));
 sky130_fd_sc_hd__a32o_2 _08350_ (.A1(_02045_),
    .A2(_02678_),
    .A3(_02777_),
    .B1(_02408_),
    .B2(_02116_),
    .X(_02778_));
 sky130_fd_sc_hd__a311o_2 _08351_ (.A1(_02523_),
    .A2(_02775_),
    .A3(_02776_),
    .B1(_02778_),
    .C1(_02454_),
    .X(_02779_));
 sky130_fd_sc_hd__o21a_2 _08352_ (.A1(_02682_),
    .A2(_02770_),
    .B1(_02779_),
    .X(_01557_));
 sky130_fd_sc_hd__and2_2 _08353_ (.A(_02532_),
    .B(\core.count_cycle[55] ),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_2 _08354_ (.A1(\core.count_instr[23] ),
    .A2(_02684_),
    .B1(_02486_),
    .B2(\core.count_instr[55] ),
    .X(_02781_));
 sky130_fd_sc_hd__a211o_2 _08355_ (.A1(\core.count_cycle[23] ),
    .A2(_02530_),
    .B1(_02780_),
    .C1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__or2_2 _08356_ (.A(\core.reg_pc[23] ),
    .B(\core.decoded_imm[23] ),
    .X(_02783_));
 sky130_fd_sc_hd__nand2_2 _08357_ (.A(\core.reg_pc[23] ),
    .B(\core.decoded_imm[23] ),
    .Y(_02784_));
 sky130_fd_sc_hd__nand2_2 _08358_ (.A(_02783_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__a21oi_2 _08359_ (.A1(_02773_),
    .A2(_02776_),
    .B1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__a31o_2 _08360_ (.A1(_02773_),
    .A2(_02776_),
    .A3(_02785_),
    .B1(_02234_),
    .X(_02787_));
 sky130_fd_sc_hd__a21oi_2 _08361_ (.A1(mem_rdata[23]),
    .A2(_02695_),
    .B1(_02675_),
    .Y(_02788_));
 sky130_fd_sc_hd__o2bb2a_2 _08362_ (.A1_N(_02546_),
    .A2_N(_02270_),
    .B1(_02707_),
    .B2(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__o211ai_2 _08363_ (.A1(_02786_),
    .A2(_02787_),
    .B1(_02789_),
    .C1(_02682_),
    .Y(_02790_));
 sky130_fd_sc_hd__o21a_2 _08364_ (.A1(_02682_),
    .A2(_02782_),
    .B1(_02790_),
    .X(_01558_));
 sky130_fd_sc_hd__nand2_2 _08365_ (.A(\core.reg_pc[24] ),
    .B(\core.decoded_imm[24] ),
    .Y(_02791_));
 sky130_fd_sc_hd__or2_2 _08366_ (.A(\core.reg_pc[24] ),
    .B(\core.decoded_imm[24] ),
    .X(_02792_));
 sky130_fd_sc_hd__and2_2 _08367_ (.A(_02791_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__or2_2 _08368_ (.A(_02774_),
    .B(_02785_),
    .X(_02794_));
 sky130_fd_sc_hd__and4b_2 _08369_ (.A_N(_02794_),
    .B(_02741_),
    .C(_02740_),
    .D(_02759_),
    .X(_02795_));
 sky130_fd_sc_hd__o21a_2 _08370_ (.A1(_02741_),
    .A2(_02758_),
    .B1(_02756_),
    .X(_02796_));
 sky130_fd_sc_hd__and3_2 _08371_ (.A(\core.reg_pc[22] ),
    .B(\core.decoded_imm[22] ),
    .C(_02783_),
    .X(_02797_));
 sky130_fd_sc_hd__a221o_2 _08372_ (.A1(\core.reg_pc[23] ),
    .A2(\core.decoded_imm[23] ),
    .B1(_02746_),
    .B2(_02795_),
    .C1(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__o21bai_2 _08373_ (.A1(_02794_),
    .A2(_02796_),
    .B1_N(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__a31o_2 _08374_ (.A1(_02690_),
    .A2(_02744_),
    .A3(_02795_),
    .B1(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_2 _08375_ (.A(_02793_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__and2_2 _08376_ (.A(\core.cpu_state[3] ),
    .B(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__o21a_2 _08377_ (.A1(_02793_),
    .A2(_02800_),
    .B1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__a21o_2 _08378_ (.A1(mem_rdata[24]),
    .A2(_02722_),
    .B1(_02709_),
    .X(_02804_));
 sky130_fd_sc_hd__a32o_2 _08379_ (.A1(_02480_),
    .A2(_02678_),
    .A3(_02804_),
    .B1(_02256_),
    .B2(_02208_),
    .X(_02805_));
 sky130_fd_sc_hd__a22o_2 _08380_ (.A1(\core.count_instr[56] ),
    .A2(_02455_),
    .B1(_02489_),
    .B2(\core.count_cycle[56] ),
    .X(_02806_));
 sky130_fd_sc_hd__a211o_2 _08381_ (.A1(\core.count_instr[24] ),
    .A2(_02684_),
    .B1(_02488_),
    .C1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__a21o_2 _08382_ (.A1(\core.count_cycle[24] ),
    .A2(_02530_),
    .B1(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__o31a_2 _08383_ (.A1(_02454_),
    .A2(_02803_),
    .A3(_02805_),
    .B1(_02808_),
    .X(_01559_));
 sky130_fd_sc_hd__and2_2 _08384_ (.A(\core.reg_pc[25] ),
    .B(\core.decoded_imm[25] ),
    .X(_02809_));
 sky130_fd_sc_hd__nor2_2 _08385_ (.A(\core.reg_pc[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_02810_));
 sky130_fd_sc_hd__or2_2 _08386_ (.A(_02809_),
    .B(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__nand2_2 _08387_ (.A(_02791_),
    .B(_02801_),
    .Y(_02812_));
 sky130_fd_sc_hd__xnor2_2 _08388_ (.A(_02811_),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__buf_1 _08389_ (.A(\core.pcpi_rs1[25] ),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_2 _08390_ (.A1(\core.count_instr[25] ),
    .A2(_02515_),
    .B1(\core.instr_rdinstrh ),
    .B2(\core.count_instr[57] ),
    .X(_02815_));
 sky130_fd_sc_hd__a221o_2 _08391_ (.A1(_02532_),
    .A2(\core.count_cycle[57] ),
    .B1(\core.count_cycle[25] ),
    .B2(_02458_),
    .C1(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__a21oi_2 _08392_ (.A1(mem_rdata[25]),
    .A2(_02708_),
    .B1(_02709_),
    .Y(_02817_));
 sky130_fd_sc_hd__nor2_2 _08393_ (.A(_02707_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__a221o_2 _08394_ (.A1(_02208_),
    .A2(_02814_),
    .B1(_02514_),
    .B2(_02816_),
    .C1(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__a21o_2 _08395_ (.A1(_02451_),
    .A2(_02813_),
    .B1(_02819_),
    .X(_01560_));
 sky130_fd_sc_hd__nor2_2 _08396_ (.A(_02809_),
    .B(_02812_),
    .Y(_02820_));
 sky130_fd_sc_hd__or2_2 _08397_ (.A(\core.reg_pc[26] ),
    .B(\core.decoded_imm[26] ),
    .X(_02821_));
 sky130_fd_sc_hd__nand2_2 _08398_ (.A(\core.reg_pc[26] ),
    .B(\core.decoded_imm[26] ),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_2 _08399_ (.A(_02821_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__o21ai_2 _08400_ (.A1(_02810_),
    .A2(_02820_),
    .B1(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__or3_2 _08401_ (.A(_02810_),
    .B(_02823_),
    .C(_02820_),
    .X(_02825_));
 sky130_fd_sc_hd__and3_2 _08402_ (.A(_02450_),
    .B(_02824_),
    .C(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__a21o_2 _08403_ (.A1(mem_rdata[26]),
    .A2(_02722_),
    .B1(_02709_),
    .X(_02827_));
 sky130_fd_sc_hd__a32o_2 _08404_ (.A1(_02480_),
    .A2(_02678_),
    .A3(_02827_),
    .B1(_02422_),
    .B2(_02208_),
    .X(_02828_));
 sky130_fd_sc_hd__a22o_2 _08405_ (.A1(\core.count_instr[26] ),
    .A2(_02515_),
    .B1(_02489_),
    .B2(\core.count_cycle[58] ),
    .X(_02829_));
 sky130_fd_sc_hd__a211o_2 _08406_ (.A1(\core.count_instr[58] ),
    .A2(_02486_),
    .B1(_02488_),
    .C1(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__a21o_2 _08407_ (.A1(\core.count_cycle[26] ),
    .A2(_02530_),
    .B1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__o31a_2 _08408_ (.A1(_02454_),
    .A2(_02826_),
    .A3(_02828_),
    .B1(_02831_),
    .X(_01561_));
 sky130_fd_sc_hd__or2_2 _08409_ (.A(\core.reg_pc[27] ),
    .B(\core.decoded_imm[27] ),
    .X(_02832_));
 sky130_fd_sc_hd__nand2_2 _08410_ (.A(\core.reg_pc[27] ),
    .B(\core.decoded_imm[27] ),
    .Y(_02833_));
 sky130_fd_sc_hd__nand2_2 _08411_ (.A(_02832_),
    .B(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__a21oi_2 _08412_ (.A1(_02822_),
    .A2(_02825_),
    .B1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__a31o_2 _08413_ (.A1(_02822_),
    .A2(_02825_),
    .A3(_02834_),
    .B1(_02234_),
    .X(_02836_));
 sky130_fd_sc_hd__or2_2 _08414_ (.A(_02835_),
    .B(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__buf_1 _08415_ (.A(\core.pcpi_rs1[27] ),
    .X(_02838_));
 sky130_fd_sc_hd__a21oi_2 _08416_ (.A1(mem_rdata[27]),
    .A2(_02708_),
    .B1(_02709_),
    .Y(_02839_));
 sky130_fd_sc_hd__o2bb2a_2 _08417_ (.A1_N(_02463_),
    .A2_N(_02838_),
    .B1(_02707_),
    .B2(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a22o_2 _08418_ (.A1(\core.count_instr[27] ),
    .A2(_02459_),
    .B1(_02489_),
    .B2(\core.count_cycle[59] ),
    .X(_02841_));
 sky130_fd_sc_hd__a211o_2 _08419_ (.A1(\core.count_instr[59] ),
    .A2(_02456_),
    .B1(_02488_),
    .C1(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__a21oi_2 _08420_ (.A1(\core.count_cycle[27] ),
    .A2(_02485_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a31oi_2 _08421_ (.A1(_02682_),
    .A2(_02837_),
    .A3(_02840_),
    .B1(_02843_),
    .Y(_01562_));
 sky130_fd_sc_hd__and2_2 _08422_ (.A(\core.count_instr[28] ),
    .B(_02684_),
    .X(_02844_));
 sky130_fd_sc_hd__a22o_2 _08423_ (.A1(\core.count_instr[60] ),
    .A2(_02486_),
    .B1(_02532_),
    .B2(\core.count_cycle[60] ),
    .X(_02845_));
 sky130_fd_sc_hd__a211o_2 _08424_ (.A1(\core.count_cycle[28] ),
    .A2(_02530_),
    .B1(_02844_),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__or3_2 _08425_ (.A(_02811_),
    .B(_02823_),
    .C(_02834_),
    .X(_02847_));
 sky130_fd_sc_hd__nor2_2 _08426_ (.A(_02823_),
    .B(_02834_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand2_2 _08427_ (.A(\core.reg_pc[25] ),
    .B(\core.decoded_imm[25] ),
    .Y(_02849_));
 sky130_fd_sc_hd__a21oi_2 _08428_ (.A1(_02791_),
    .A2(_02849_),
    .B1(_02810_),
    .Y(_02850_));
 sky130_fd_sc_hd__and3_2 _08429_ (.A(\core.reg_pc[26] ),
    .B(\core.decoded_imm[26] ),
    .C(_02832_),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_2 _08430_ (.A1(\core.reg_pc[27] ),
    .A2(\core.decoded_imm[27] ),
    .B1(_02848_),
    .B2(_02850_),
    .C1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__o21bai_2 _08431_ (.A1(_02801_),
    .A2(_02847_),
    .B1_N(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__nor2_2 _08432_ (.A(\core.reg_pc[28] ),
    .B(\core.decoded_imm[28] ),
    .Y(_02854_));
 sky130_fd_sc_hd__and2_2 _08433_ (.A(\core.reg_pc[28] ),
    .B(\core.decoded_imm[28] ),
    .X(_02855_));
 sky130_fd_sc_hd__nor2_2 _08434_ (.A(_02854_),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__or2_2 _08435_ (.A(_02853_),
    .B(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__nand2_2 _08436_ (.A(_02853_),
    .B(_02856_),
    .Y(_02858_));
 sky130_fd_sc_hd__a21o_2 _08437_ (.A1(mem_rdata[28]),
    .A2(_02464_),
    .B1(_02675_),
    .X(_02859_));
 sky130_fd_sc_hd__a32o_2 _08438_ (.A1(_02045_),
    .A2(_02678_),
    .A3(_02859_),
    .B1(_02246_),
    .B2(_02116_),
    .X(_02860_));
 sky130_fd_sc_hd__a311o_2 _08439_ (.A1(_02523_),
    .A2(_02857_),
    .A3(_02858_),
    .B1(_02860_),
    .C1(_02454_),
    .X(_02861_));
 sky130_fd_sc_hd__o21a_2 _08440_ (.A1(_02682_),
    .A2(_02846_),
    .B1(_02861_),
    .X(_01563_));
 sky130_fd_sc_hd__and2_2 _08441_ (.A(\core.count_instr[61] ),
    .B(_02486_),
    .X(_02862_));
 sky130_fd_sc_hd__a22o_2 _08442_ (.A1(\core.count_instr[29] ),
    .A2(_02684_),
    .B1(_02532_),
    .B2(\core.count_cycle[61] ),
    .X(_02863_));
 sky130_fd_sc_hd__a211o_2 _08443_ (.A1(\core.count_cycle[29] ),
    .A2(_02530_),
    .B1(_02862_),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__or2_2 _08444_ (.A(\core.reg_pc[29] ),
    .B(\core.decoded_imm[29] ),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_2 _08445_ (.A(\core.reg_pc[29] ),
    .B(\core.decoded_imm[29] ),
    .Y(_02866_));
 sky130_fd_sc_hd__a21o_2 _08446_ (.A1(_02853_),
    .A2(_02856_),
    .B1(_02855_),
    .X(_02867_));
 sky130_fd_sc_hd__a21oi_2 _08447_ (.A1(_02865_),
    .A2(_02866_),
    .B1(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__a31o_2 _08448_ (.A1(_02865_),
    .A2(_02866_),
    .A3(_02867_),
    .B1(_02234_),
    .X(_02869_));
 sky130_fd_sc_hd__a21oi_2 _08449_ (.A1(mem_rdata[29]),
    .A2(_02695_),
    .B1(_02675_),
    .Y(_02870_));
 sky130_fd_sc_hd__o2bb2a_2 _08450_ (.A1_N(_02546_),
    .A2_N(_02414_),
    .B1(_02707_),
    .B2(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__o211ai_2 _08451_ (.A1(_02868_),
    .A2(_02869_),
    .B1(_02871_),
    .C1(_02531_),
    .Y(_02872_));
 sky130_fd_sc_hd__o21a_2 _08452_ (.A1(_02682_),
    .A2(_02864_),
    .B1(_02872_),
    .X(_01564_));
 sky130_fd_sc_hd__and2_2 _08453_ (.A(\core.count_instr[62] ),
    .B(_02486_),
    .X(_02873_));
 sky130_fd_sc_hd__a22o_2 _08454_ (.A1(\core.count_instr[30] ),
    .A2(_02684_),
    .B1(_02532_),
    .B2(\core.count_cycle[62] ),
    .X(_02874_));
 sky130_fd_sc_hd__a211o_2 _08455_ (.A1(\core.count_cycle[30] ),
    .A2(_02458_),
    .B1(_02873_),
    .C1(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__nand2_2 _08456_ (.A(\core.reg_pc[30] ),
    .B(\core.decoded_imm[30] ),
    .Y(_02876_));
 sky130_fd_sc_hd__or2_2 _08457_ (.A(\core.reg_pc[30] ),
    .B(\core.decoded_imm[30] ),
    .X(_02877_));
 sky130_fd_sc_hd__nand2_2 _08458_ (.A(_02876_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_2 _08459_ (.A(_02865_),
    .B(_02867_),
    .Y(_02879_));
 sky130_fd_sc_hd__and3_2 _08460_ (.A(_02866_),
    .B(_02878_),
    .C(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__a21o_2 _08461_ (.A1(_02866_),
    .A2(_02879_),
    .B1(_02878_),
    .X(_02881_));
 sky130_fd_sc_hd__nand2_2 _08462_ (.A(_02523_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__a21oi_2 _08463_ (.A1(mem_rdata[30]),
    .A2(_02695_),
    .B1(_02675_),
    .Y(_02883_));
 sky130_fd_sc_hd__o2bb2a_2 _08464_ (.A1_N(_02546_),
    .A2_N(_02242_),
    .B1(_02707_),
    .B2(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__o211ai_2 _08465_ (.A1(_02880_),
    .A2(_02882_),
    .B1(_02884_),
    .C1(_02531_),
    .Y(_02885_));
 sky130_fd_sc_hd__o21a_2 _08466_ (.A1(_02682_),
    .A2(_02875_),
    .B1(_02885_),
    .X(_01566_));
 sky130_fd_sc_hd__xnor2_2 _08467_ (.A(\core.reg_pc[31] ),
    .B(\core.decoded_imm[31] ),
    .Y(_02886_));
 sky130_fd_sc_hd__a21oi_2 _08468_ (.A1(_02876_),
    .A2(_02881_),
    .B1(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__a31o_2 _08469_ (.A1(_02876_),
    .A2(_02881_),
    .A3(_02886_),
    .B1(_02234_),
    .X(_02888_));
 sky130_fd_sc_hd__and2_2 _08470_ (.A(\core.count_instr[63] ),
    .B(\core.instr_rdinstrh ),
    .X(_02889_));
 sky130_fd_sc_hd__a22o_2 _08471_ (.A1(\core.count_instr[31] ),
    .A2(_02515_),
    .B1(_02489_),
    .B2(\core.count_cycle[63] ),
    .X(_02890_));
 sky130_fd_sc_hd__a211o_2 _08472_ (.A1(\core.count_cycle[31] ),
    .A2(_02458_),
    .B1(_02889_),
    .C1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__a21oi_2 _08473_ (.A1(mem_rdata[31]),
    .A2(_02722_),
    .B1(_02709_),
    .Y(_02892_));
 sky130_fd_sc_hd__nor2_2 _08474_ (.A(_02707_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__a221o_2 _08475_ (.A1(_02208_),
    .A2(_02237_),
    .B1(_02514_),
    .B2(_02891_),
    .C1(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__o21bai_2 _08476_ (.A1(_02887_),
    .A2(_02888_),
    .B1_N(_02894_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2_2 _08477_ (.A(\core.instr_or ),
    .B(\core.instr_ori ),
    .X(_02895_));
 sky130_fd_sc_hd__or2_2 _08478_ (.A(\core.instr_xori ),
    .B(\core.instr_xor ),
    .X(_02896_));
 sky130_fd_sc_hd__or2_2 _08479_ (.A(\core.instr_andi ),
    .B(\core.instr_and ),
    .X(_02897_));
 sky130_fd_sc_hd__buf_1 _08480_ (.A(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__nor4_2 _08481_ (.A(\core.is_compare ),
    .B(_02895_),
    .C(_02896_),
    .D(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__buf_1 _08482_ (.A(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__buf_1 _08483_ (.A(_02895_),
    .X(_02901_));
 sky130_fd_sc_hd__buf_1 _08484_ (.A(_02896_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_2 _08485_ (.A0(_02898_),
    .A1(_02902_),
    .S(_02434_),
    .X(_02903_));
 sky130_fd_sc_hd__o21a_2 _08486_ (.A1(_02901_),
    .A2(_02903_),
    .B1(_02435_),
    .X(_02904_));
 sky130_fd_sc_hd__a221o_2 _08487_ (.A1(\core.is_compare ),
    .A2(_02445_),
    .B1(_02900_),
    .B2(_02436_),
    .C1(_02904_),
    .X(\core.alu_out[0] ));
 sky130_fd_sc_hd__buf_1 _08488_ (.A(_02898_),
    .X(_02905_));
 sky130_fd_sc_hd__buf_1 _08489_ (.A(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__nor2_2 _08490_ (.A(\core.instr_xori ),
    .B(\core.instr_xor ),
    .Y(_02907_));
 sky130_fd_sc_hd__a21oi_2 _08491_ (.A1(_02476_),
    .A2(_02366_),
    .B1(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__o22a_2 _08492_ (.A1(_02476_),
    .A2(_02366_),
    .B1(_02895_),
    .B2(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__a31o_2 _08493_ (.A1(_02476_),
    .A2(_02366_),
    .A3(_02906_),
    .B1(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__inv_2 _08494_ (.A(\core.instr_sub ),
    .Y(_02911_));
 sky130_fd_sc_hd__buf_1 _08495_ (.A(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__and3_2 _08496_ (.A(_02367_),
    .B(_02368_),
    .C(_02369_),
    .X(_02913_));
 sky130_fd_sc_hd__or2_2 _08497_ (.A(_02370_),
    .B(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__a21oi_2 _08498_ (.A1(_02912_),
    .A2(_02368_),
    .B1(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__or4_2 _08499_ (.A(\core.is_compare ),
    .B(_02895_),
    .C(_02896_),
    .D(_02897_),
    .X(_02916_));
 sky130_fd_sc_hd__buf_1 _08500_ (.A(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__a31o_2 _08501_ (.A1(_02912_),
    .A2(_02368_),
    .A3(_02914_),
    .B1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__o22a_2 _08502_ (.A1(_02900_),
    .A2(_02910_),
    .B1(_02915_),
    .B2(_02918_),
    .X(\core.alu_out[1] ));
 sky130_fd_sc_hd__a22o_2 _08503_ (.A1(\core.pcpi_rs1[0] ),
    .A2(\core.mem_la_wdata[0] ),
    .B1(\core.mem_la_wdata[1] ),
    .B2(\core.pcpi_rs1[1] ),
    .X(_02919_));
 sky130_fd_sc_hd__o21ai_2 _08504_ (.A1(\core.pcpi_rs1[1] ),
    .A2(_02366_),
    .B1(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__buf_1 _08505_ (.A(_02911_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_2 _08506_ (.A0(_02371_),
    .A1(_02920_),
    .S(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__xnor2_2 _08507_ (.A(_02364_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__buf_1 _08508_ (.A(_02896_),
    .X(_02924_));
 sky130_fd_sc_hd__a21o_2 _08509_ (.A1(_02362_),
    .A2(_02924_),
    .B1(_02901_),
    .X(_02925_));
 sky130_fd_sc_hd__a31o_2 _08510_ (.A1(\core.mem_la_wdata[2] ),
    .A2(_02372_),
    .A3(_02905_),
    .B1(_02899_),
    .X(_02926_));
 sky130_fd_sc_hd__a21oi_2 _08511_ (.A1(_02363_),
    .A2(_02925_),
    .B1(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21oi_2 _08512_ (.A1(_02900_),
    .A2(_02923_),
    .B1(_02927_),
    .Y(\core.alu_out[2] ));
 sky130_fd_sc_hd__a21bo_2 _08513_ (.A1(_02362_),
    .A2(_02920_),
    .B1_N(_02363_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_2 _08514_ (.A0(_02374_),
    .A1(_02928_),
    .S(_02921_),
    .X(_02929_));
 sky130_fd_sc_hd__xnor2_2 _08515_ (.A(_02361_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__a21o_2 _08516_ (.A1(_02359_),
    .A2(_02924_),
    .B1(_02901_),
    .X(_02931_));
 sky130_fd_sc_hd__a31o_2 _08517_ (.A1(\core.mem_la_wdata[3] ),
    .A2(_02375_),
    .A3(_02905_),
    .B1(_02899_),
    .X(_02932_));
 sky130_fd_sc_hd__a21oi_2 _08518_ (.A1(_02360_),
    .A2(_02931_),
    .B1(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__a21oi_2 _08519_ (.A1(_02900_),
    .A2(_02930_),
    .B1(_02933_),
    .Y(\core.alu_out[3] ));
 sky130_fd_sc_hd__a21bo_2 _08520_ (.A1(_02359_),
    .A2(_02928_),
    .B1_N(_02360_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_2 _08521_ (.A0(_02377_),
    .A1(_02934_),
    .S(_02921_),
    .X(_02935_));
 sky130_fd_sc_hd__xor2_2 _08522_ (.A(_02358_),
    .B(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__buf_1 _08523_ (.A(_02895_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_2 _08524_ (.A0(_02902_),
    .A1(_02897_),
    .S(_02356_),
    .X(_02938_));
 sky130_fd_sc_hd__o21ba_2 _08525_ (.A1(_02937_),
    .A2(_02938_),
    .B1_N(_02357_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_2 _08526_ (.A0(_02936_),
    .A1(_02939_),
    .S(_02917_),
    .X(_02940_));
 sky130_fd_sc_hd__buf_1 _08527_ (.A(_02940_),
    .X(\core.alu_out[4] ));
 sky130_fd_sc_hd__buf_1 _08528_ (.A(_02917_),
    .X(_02941_));
 sky130_fd_sc_hd__buf_1 _08529_ (.A(\core.instr_sub ),
    .X(_02942_));
 sky130_fd_sc_hd__nand2_2 _08530_ (.A(_02387_),
    .B(_02355_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand2_2 _08531_ (.A(_02358_),
    .B(_02377_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_2 _08532_ (.A(\core.mem_la_wdata[4] ),
    .B(\core.pcpi_rs1[4] ),
    .Y(_02945_));
 sky130_fd_sc_hd__a21o_2 _08533_ (.A1(_02945_),
    .A2(_02934_),
    .B1(_02357_),
    .X(_02946_));
 sky130_fd_sc_hd__nor2_2 _08534_ (.A(_02942_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__a31o_2 _08535_ (.A1(_02942_),
    .A2(_02943_),
    .A3(_02944_),
    .B1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__xnor2_2 _08536_ (.A(_02354_),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__buf_1 _08537_ (.A(_02937_),
    .X(_02950_));
 sky130_fd_sc_hd__a21oi_2 _08538_ (.A1(_02353_),
    .A2(_02924_),
    .B1(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__nor2_2 _08539_ (.A(_02352_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__buf_1 _08540_ (.A(_02899_),
    .X(_02953_));
 sky130_fd_sc_hd__a31o_2 _08541_ (.A1(\core.mem_la_wdata[5] ),
    .A2(_02388_),
    .A3(_02906_),
    .B1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__o22a_2 _08542_ (.A1(_02941_),
    .A2(_02949_),
    .B1(_02952_),
    .B2(_02954_),
    .X(\core.alu_out[5] ));
 sky130_fd_sc_hd__nor2_2 _08543_ (.A(_02378_),
    .B(_02390_),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ai_2 _08544_ (.A1(_02352_),
    .A2(_02946_),
    .B1(_02353_),
    .Y(_02956_));
 sky130_fd_sc_hd__mux2_2 _08545_ (.A0(_02955_),
    .A1(_02956_),
    .S(_02921_),
    .X(_02957_));
 sky130_fd_sc_hd__nor2_2 _08546_ (.A(_02386_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21o_2 _08547_ (.A1(_02386_),
    .A2(_02957_),
    .B1(_02917_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_2 _08548_ (.A0(_02905_),
    .A1(_02924_),
    .S(_02384_),
    .X(_02960_));
 sky130_fd_sc_hd__o21a_2 _08549_ (.A1(_02950_),
    .A2(_02960_),
    .B1(_02385_),
    .X(_02961_));
 sky130_fd_sc_hd__o22a_2 _08550_ (.A1(_02958_),
    .A2(_02959_),
    .B1(_02961_),
    .B2(_02900_),
    .X(\core.alu_out[6] ));
 sky130_fd_sc_hd__o21ba_2 _08551_ (.A1(_02379_),
    .A2(_02907_),
    .B1_N(_02901_),
    .X(_02962_));
 sky130_fd_sc_hd__nor2_2 _08552_ (.A(_02381_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21o_2 _08553_ (.A1(_02379_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_02964_));
 sky130_fd_sc_hd__inv_2 _08554_ (.A(_02386_),
    .Y(_02965_));
 sky130_fd_sc_hd__nor2_2 _08555_ (.A(_02965_),
    .B(_02955_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_2 _08556_ (.A(_02385_),
    .B(_02956_),
    .Y(_02967_));
 sky130_fd_sc_hd__a21o_2 _08557_ (.A1(_02384_),
    .A2(_02967_),
    .B1(\core.instr_sub ),
    .X(_02968_));
 sky130_fd_sc_hd__o31ai_2 _08558_ (.A1(_02912_),
    .A2(_02391_),
    .A3(_02966_),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xnor2_2 _08559_ (.A(_02382_),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__o22a_2 _08560_ (.A1(_02963_),
    .A2(_02964_),
    .B1(_02970_),
    .B2(_02941_),
    .X(\core.alu_out[7] ));
 sky130_fd_sc_hd__inv_2 _08561_ (.A(_02395_),
    .Y(_02971_));
 sky130_fd_sc_hd__inv_2 _08562_ (.A(_02382_),
    .Y(_02972_));
 sky130_fd_sc_hd__o211a_2 _08563_ (.A1(\core.mem_la_wdata[7] ),
    .A2(_02380_),
    .B1(\core.mem_la_wdata[6] ),
    .C1(_02383_),
    .X(_02973_));
 sky130_fd_sc_hd__a311o_2 _08564_ (.A1(_02972_),
    .A2(_02965_),
    .A3(_02956_),
    .B1(_02973_),
    .C1(_02379_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_2 _08565_ (.A0(_02971_),
    .A1(_02974_),
    .S(_02911_),
    .X(_02975_));
 sky130_fd_sc_hd__xnor2_2 _08566_ (.A(_02348_),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__mux2_2 _08567_ (.A0(_02898_),
    .A1(_02902_),
    .S(_02347_),
    .X(_02977_));
 sky130_fd_sc_hd__o21a_2 _08568_ (.A1(_02901_),
    .A2(_02977_),
    .B1(_02346_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_1 _08569_ (.A(_02916_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_2 _08570_ (.A0(_02976_),
    .A1(_02978_),
    .S(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__buf_1 _08571_ (.A(_02980_),
    .X(\core.alu_out[8] ));
 sky130_fd_sc_hd__a21oi_2 _08572_ (.A1(_02329_),
    .A2(_02924_),
    .B1(_02950_),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2_2 _08573_ (.A(_02328_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__a31o_2 _08574_ (.A1(\core.pcpi_rs2[9] ),
    .A2(_02331_),
    .A3(_02905_),
    .B1(_02953_),
    .X(_02983_));
 sky130_fd_sc_hd__and2_2 _08575_ (.A(_02348_),
    .B(_02395_),
    .X(_02984_));
 sky130_fd_sc_hd__a21o_2 _08576_ (.A1(_02326_),
    .A2(_02327_),
    .B1(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__a21boi_2 _08577_ (.A1(_02346_),
    .A2(_02974_),
    .B1_N(_02347_),
    .Y(_02986_));
 sky130_fd_sc_hd__mux2_2 _08578_ (.A0(_02985_),
    .A1(_02986_),
    .S(_02912_),
    .X(_02987_));
 sky130_fd_sc_hd__xor2_2 _08579_ (.A(_02330_),
    .B(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__o22a_2 _08580_ (.A1(_02982_),
    .A2(_02983_),
    .B1(_02988_),
    .B2(_02941_),
    .X(\core.alu_out[9] ));
 sky130_fd_sc_hd__a21o_2 _08581_ (.A1(_02330_),
    .A2(_02985_),
    .B1(_02332_),
    .X(_02989_));
 sky130_fd_sc_hd__inv_2 _08582_ (.A(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__a21oi_2 _08583_ (.A1(_02329_),
    .A2(_02986_),
    .B1(_02328_),
    .Y(_02991_));
 sky130_fd_sc_hd__mux2_2 _08584_ (.A0(_02990_),
    .A1(_02991_),
    .S(_02911_),
    .X(_02992_));
 sky130_fd_sc_hd__xnor2_2 _08585_ (.A(_02325_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__and2_2 _08586_ (.A(\core.pcpi_rs2[10] ),
    .B(_02323_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_2 _08587_ (.A0(_02902_),
    .A1(_02898_),
    .S(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__o21a_2 _08588_ (.A1(_02901_),
    .A2(_02995_),
    .B1(_02322_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_2 _08589_ (.A0(_02993_),
    .A1(_02996_),
    .S(_02979_),
    .X(_02997_));
 sky130_fd_sc_hd__buf_1 _08590_ (.A(_02997_),
    .X(\core.alu_out[10] ));
 sky130_fd_sc_hd__nor2_2 _08591_ (.A(_02319_),
    .B(_02907_),
    .Y(_02998_));
 sky130_fd_sc_hd__o21ba_2 _08592_ (.A1(_02950_),
    .A2(_02998_),
    .B1_N(_02320_),
    .X(_02999_));
 sky130_fd_sc_hd__a21o_2 _08593_ (.A1(_02319_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_03000_));
 sky130_fd_sc_hd__o21ai_2 _08594_ (.A1(_02994_),
    .A2(_02991_),
    .B1(_02322_),
    .Y(_03001_));
 sky130_fd_sc_hd__a21o_2 _08595_ (.A1(_02325_),
    .A2(_02989_),
    .B1(_02334_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_2 _08596_ (.A0(_03001_),
    .A1(_03002_),
    .S(_02942_),
    .X(_03003_));
 sky130_fd_sc_hd__xor2_2 _08597_ (.A(_02321_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__o22a_2 _08598_ (.A1(_02999_),
    .A2(_03000_),
    .B1(_03004_),
    .B2(_02941_),
    .X(\core.alu_out[11] ));
 sky130_fd_sc_hd__or4_2 _08599_ (.A(_02321_),
    .B(_02325_),
    .C(_02330_),
    .D(_02348_),
    .X(_03005_));
 sky130_fd_sc_hd__inv_2 _08600_ (.A(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__o21ai_2 _08601_ (.A1(_02328_),
    .A2(_02347_),
    .B1(_02329_),
    .Y(_03007_));
 sky130_fd_sc_hd__o221a_2 _08602_ (.A1(\core.pcpi_rs2[11] ),
    .A2(_02336_),
    .B1(_02994_),
    .B2(_03007_),
    .C1(_02322_),
    .X(_03008_));
 sky130_fd_sc_hd__a211oi_2 _08603_ (.A1(_02974_),
    .A2(_03006_),
    .B1(_03008_),
    .C1(_02319_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21o_2 _08604_ (.A1(_02321_),
    .A2(_03002_),
    .B1(_02337_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_2 _08605_ (.A0(_03009_),
    .A1(_03010_),
    .S(\core.instr_sub ),
    .X(_03011_));
 sky130_fd_sc_hd__xor2_2 _08606_ (.A(_02318_),
    .B(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_2 _08607_ (.A0(_02898_),
    .A1(_02896_),
    .S(_02317_),
    .X(_03013_));
 sky130_fd_sc_hd__o21ba_2 _08608_ (.A1(_02937_),
    .A2(_03013_),
    .B1_N(_02316_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_2 _08609_ (.A0(_03012_),
    .A1(_03014_),
    .S(_02979_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_1 _08610_ (.A(_03015_),
    .X(\core.alu_out[12] ));
 sky130_fd_sc_hd__a21oi_2 _08611_ (.A1(_02313_),
    .A2(_02924_),
    .B1(_02950_),
    .Y(_03016_));
 sky130_fd_sc_hd__nor2_2 _08612_ (.A(_02311_),
    .B(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__a31o_2 _08613_ (.A1(\core.pcpi_rs2[13] ),
    .A2(_02312_),
    .A3(_02905_),
    .B1(_02953_),
    .X(_03018_));
 sky130_fd_sc_hd__and2_2 _08614_ (.A(_02318_),
    .B(_03010_),
    .X(_03019_));
 sky130_fd_sc_hd__a21o_2 _08615_ (.A1(_02339_),
    .A2(_02315_),
    .B1(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__o21a_2 _08616_ (.A1(_02316_),
    .A2(_03009_),
    .B1(_02317_),
    .X(_03021_));
 sky130_fd_sc_hd__mux2_2 _08617_ (.A0(_03020_),
    .A1(_03021_),
    .S(_02912_),
    .X(_03022_));
 sky130_fd_sc_hd__xor2_2 _08618_ (.A(_02314_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__o22a_2 _08619_ (.A1(_03017_),
    .A2(_03018_),
    .B1(_03023_),
    .B2(_02941_),
    .X(\core.alu_out[13] ));
 sky130_fd_sc_hd__a21oi_2 _08620_ (.A1(_02314_),
    .A2(_03020_),
    .B1(_02340_),
    .Y(_03024_));
 sky130_fd_sc_hd__o21a_2 _08621_ (.A1(_02311_),
    .A2(_03021_),
    .B1(_02313_),
    .X(_03025_));
 sky130_fd_sc_hd__inv_2 _08622_ (.A(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__mux2_2 _08623_ (.A0(_03024_),
    .A1(_03026_),
    .S(_02911_),
    .X(_03027_));
 sky130_fd_sc_hd__xnor2_2 _08624_ (.A(_02310_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__mux2_2 _08625_ (.A0(_02898_),
    .A1(_02902_),
    .S(_02307_),
    .X(_03029_));
 sky130_fd_sc_hd__o21a_2 _08626_ (.A1(_02937_),
    .A2(_03029_),
    .B1(_02309_),
    .X(_03030_));
 sky130_fd_sc_hd__mux2_2 _08627_ (.A0(_03028_),
    .A1(_03030_),
    .S(_02979_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_1 _08628_ (.A(_03031_),
    .X(\core.alu_out[14] ));
 sky130_fd_sc_hd__a21oi_2 _08629_ (.A1(_02307_),
    .A2(_02309_),
    .B1(_03024_),
    .Y(_03032_));
 sky130_fd_sc_hd__a211o_2 _08630_ (.A1(_02307_),
    .A2(_03025_),
    .B1(_02308_),
    .C1(\core.instr_sub ),
    .X(_03033_));
 sky130_fd_sc_hd__o31a_2 _08631_ (.A1(_02912_),
    .A2(_02343_),
    .A3(_03032_),
    .B1(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__xor2_2 _08632_ (.A(_02305_),
    .B(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__o21ba_2 _08633_ (.A1(_02303_),
    .A2(_02907_),
    .B1_N(_02901_),
    .X(_03036_));
 sky130_fd_sc_hd__nor2_2 _08634_ (.A(_02304_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__a21o_2 _08635_ (.A1(_02303_),
    .A2(_02906_),
    .B1(_02900_),
    .X(_03038_));
 sky130_fd_sc_hd__o22a_2 _08636_ (.A1(_02941_),
    .A2(_03035_),
    .B1(_03037_),
    .B2(_03038_),
    .X(\core.alu_out[15] ));
 sky130_fd_sc_hd__inv_2 _08637_ (.A(_02397_),
    .Y(_03039_));
 sky130_fd_sc_hd__or4_2 _08638_ (.A(_02305_),
    .B(_02310_),
    .C(_02314_),
    .D(_02318_),
    .X(_03040_));
 sky130_fd_sc_hd__o211a_2 _08639_ (.A1(_02311_),
    .A2(_02317_),
    .B1(_02313_),
    .C1(_02307_),
    .X(_03041_));
 sky130_fd_sc_hd__or3_2 _08640_ (.A(_02304_),
    .B(_02308_),
    .C(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__o221a_2 _08641_ (.A1(_02301_),
    .A2(_02302_),
    .B1(_03009_),
    .B2(_03040_),
    .C1(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__mux2_2 _08642_ (.A0(_03039_),
    .A1(_03043_),
    .S(_02911_),
    .X(_03044_));
 sky130_fd_sc_hd__xnor2_2 _08643_ (.A(_02400_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__mux2_2 _08644_ (.A0(_02902_),
    .A1(_02897_),
    .S(_02399_),
    .X(_03046_));
 sky130_fd_sc_hd__o21ba_2 _08645_ (.A1(_02937_),
    .A2(_03046_),
    .B1_N(_02398_),
    .X(_03047_));
 sky130_fd_sc_hd__mux2_2 _08646_ (.A0(_03045_),
    .A1(_03047_),
    .S(_02979_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_1 _08647_ (.A(_03048_),
    .X(\core.alu_out[16] ));
 sky130_fd_sc_hd__and2_2 _08648_ (.A(\core.pcpi_rs2[17] ),
    .B(_02293_),
    .X(_03049_));
 sky130_fd_sc_hd__nor2_2 _08649_ (.A(_03049_),
    .B(_02907_),
    .Y(_03050_));
 sky130_fd_sc_hd__o21a_2 _08650_ (.A1(_02950_),
    .A2(_03050_),
    .B1(_02292_),
    .X(_03051_));
 sky130_fd_sc_hd__a21o_2 _08651_ (.A1(_03049_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_03052_));
 sky130_fd_sc_hd__a2bb2o_2 _08652_ (.A1_N(_02397_),
    .A2_N(_02400_),
    .B1(_02290_),
    .B2(_02291_),
    .X(_03053_));
 sky130_fd_sc_hd__inv_2 _08653_ (.A(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__o21bai_2 _08654_ (.A1(_02398_),
    .A2(_03043_),
    .B1_N(_02399_),
    .Y(_03055_));
 sky130_fd_sc_hd__mux2_2 _08655_ (.A0(_03054_),
    .A1(_03055_),
    .S(_02921_),
    .X(_03056_));
 sky130_fd_sc_hd__xnor2_2 _08656_ (.A(_02295_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__o22a_2 _08657_ (.A1(_03051_),
    .A2(_03052_),
    .B1(_03057_),
    .B2(_02941_),
    .X(\core.alu_out[17] ));
 sky130_fd_sc_hd__a21o_2 _08658_ (.A1(_02295_),
    .A2(_03053_),
    .B1(_02296_),
    .X(_03058_));
 sky130_fd_sc_hd__o21ai_2 _08659_ (.A1(_03049_),
    .A2(_03055_),
    .B1(_02292_),
    .Y(_03059_));
 sky130_fd_sc_hd__mux2_2 _08660_ (.A0(_03058_),
    .A1(_03059_),
    .S(_02921_),
    .X(_03060_));
 sky130_fd_sc_hd__xor2_2 _08661_ (.A(_02289_),
    .B(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_2 _08662_ (.A0(_02897_),
    .A1(_02896_),
    .S(_02288_),
    .X(_03062_));
 sky130_fd_sc_hd__o21ba_2 _08663_ (.A1(_02937_),
    .A2(_03062_),
    .B1_N(_02287_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_2 _08664_ (.A0(_03061_),
    .A1(_03063_),
    .S(_02979_),
    .X(_03064_));
 sky130_fd_sc_hd__buf_1 _08665_ (.A(_03064_),
    .X(\core.alu_out[18] ));
 sky130_fd_sc_hd__a21oi_2 _08666_ (.A1(\core.pcpi_rs2[19] ),
    .A2(_02736_),
    .B1(_02907_),
    .Y(_03065_));
 sky130_fd_sc_hd__o22a_2 _08667_ (.A1(\core.pcpi_rs2[19] ),
    .A2(_02736_),
    .B1(_02895_),
    .B2(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__a31o_2 _08668_ (.A1(\core.pcpi_rs2[19] ),
    .A2(_02736_),
    .A3(_02905_),
    .B1(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__a211o_2 _08669_ (.A1(_02289_),
    .A2(_03058_),
    .B1(_02912_),
    .C1(_02299_),
    .X(_03068_));
 sky130_fd_sc_hd__a211o_2 _08670_ (.A1(_02288_),
    .A2(_03059_),
    .B1(_02942_),
    .C1(_02287_),
    .X(_03069_));
 sky130_fd_sc_hd__a21oi_2 _08671_ (.A1(_03068_),
    .A2(_03069_),
    .B1(_02286_),
    .Y(_03070_));
 sky130_fd_sc_hd__a31o_2 _08672_ (.A1(_02286_),
    .A2(_03068_),
    .A3(_03069_),
    .B1(_02917_),
    .X(_03071_));
 sky130_fd_sc_hd__o22a_2 _08673_ (.A1(_02900_),
    .A2(_03067_),
    .B1(_03070_),
    .B2(_03071_),
    .X(\core.alu_out[19] ));
 sky130_fd_sc_hd__inv_2 _08674_ (.A(_02404_),
    .Y(_03072_));
 sky130_fd_sc_hd__a221o_2 _08675_ (.A1(\core.pcpi_rs2[18] ),
    .A2(_02298_),
    .B1(_02292_),
    .B2(_02399_),
    .C1(_03049_),
    .X(_03073_));
 sky130_fd_sc_hd__o221a_2 _08676_ (.A1(\core.pcpi_rs2[19] ),
    .A2(\core.pcpi_rs1[19] ),
    .B1(\core.pcpi_rs2[18] ),
    .B2(_02298_),
    .C1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__a21oi_2 _08677_ (.A1(\core.pcpi_rs2[19] ),
    .A2(\core.pcpi_rs1[19] ),
    .B1(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__or3b_2 _08678_ (.A(_02289_),
    .B(_02295_),
    .C_N(_02400_),
    .X(_03076_));
 sky130_fd_sc_hd__or3b_2 _08679_ (.A(_03043_),
    .B(_03076_),
    .C_N(_02286_),
    .X(_03077_));
 sky130_fd_sc_hd__nand2_2 _08680_ (.A(_03075_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__mux2_2 _08681_ (.A0(_03072_),
    .A1(_03078_),
    .S(_02911_),
    .X(_03079_));
 sky130_fd_sc_hd__xnor2_2 _08682_ (.A(_02279_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__mux2_2 _08683_ (.A0(_02898_),
    .A1(_02902_),
    .S(_02278_),
    .X(_03081_));
 sky130_fd_sc_hd__o21a_2 _08684_ (.A1(_02937_),
    .A2(_03081_),
    .B1(_02276_),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_2 _08685_ (.A0(_03080_),
    .A1(_03082_),
    .S(_02979_),
    .X(_03083_));
 sky130_fd_sc_hd__buf_1 _08686_ (.A(_03083_),
    .X(\core.alu_out[20] ));
 sky130_fd_sc_hd__a21oi_2 _08687_ (.A1(_02282_),
    .A2(_02924_),
    .B1(_02901_),
    .Y(_03084_));
 sky130_fd_sc_hd__nor2_2 _08688_ (.A(_02280_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__a31o_2 _08689_ (.A1(\core.pcpi_rs2[21] ),
    .A2(_02281_),
    .A3(_02905_),
    .B1(_02953_),
    .X(_03086_));
 sky130_fd_sc_hd__and2_2 _08690_ (.A(_02279_),
    .B(_02404_),
    .X(_03087_));
 sky130_fd_sc_hd__a21o_2 _08691_ (.A1(_02405_),
    .A2(_02277_),
    .B1(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a21boi_2 _08692_ (.A1(_02276_),
    .A2(_03078_),
    .B1_N(_02278_),
    .Y(_03089_));
 sky130_fd_sc_hd__mux2_2 _08693_ (.A0(_03088_),
    .A1(_03089_),
    .S(_02912_),
    .X(_03090_));
 sky130_fd_sc_hd__xor2_2 _08694_ (.A(_02283_),
    .B(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__o22a_2 _08695_ (.A1(_03085_),
    .A2(_03086_),
    .B1(_03091_),
    .B2(_02941_),
    .X(\core.alu_out[21] ));
 sky130_fd_sc_hd__a21oi_2 _08696_ (.A1(_02283_),
    .A2(_03088_),
    .B1(_02406_),
    .Y(_03092_));
 sky130_fd_sc_hd__o21ai_2 _08697_ (.A1(_02280_),
    .A2(_03089_),
    .B1(_02282_),
    .Y(_03093_));
 sky130_fd_sc_hd__mux2_2 _08698_ (.A0(_03092_),
    .A1(_03093_),
    .S(_02921_),
    .X(_03094_));
 sky130_fd_sc_hd__nor2_2 _08699_ (.A(_02275_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a21o_2 _08700_ (.A1(_02275_),
    .A2(_03094_),
    .B1(_02917_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_2 _08701_ (.A0(_02902_),
    .A1(_02898_),
    .S(_02273_),
    .X(_03097_));
 sky130_fd_sc_hd__o21ba_2 _08702_ (.A1(_02950_),
    .A2(_03097_),
    .B1_N(_02274_),
    .X(_03098_));
 sky130_fd_sc_hd__o22a_2 _08703_ (.A1(_03095_),
    .A2(_03096_),
    .B1(_03098_),
    .B2(_02900_),
    .X(\core.alu_out[22] ));
 sky130_fd_sc_hd__nor2_2 _08704_ (.A(_02273_),
    .B(_03093_),
    .Y(_03099_));
 sky130_fd_sc_hd__inv_2 _08705_ (.A(_03092_),
    .Y(_03100_));
 sky130_fd_sc_hd__a211o_2 _08706_ (.A1(_02275_),
    .A2(_03100_),
    .B1(_02409_),
    .C1(_02921_),
    .X(_03101_));
 sky130_fd_sc_hd__o31a_2 _08707_ (.A1(_02942_),
    .A2(_02274_),
    .A3(_03099_),
    .B1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__xor2_2 _08708_ (.A(_02272_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__o21ba_2 _08709_ (.A1(_02269_),
    .A2(_02907_),
    .B1_N(_02901_),
    .X(_03104_));
 sky130_fd_sc_hd__nor2_2 _08710_ (.A(_02271_),
    .B(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__a21o_2 _08711_ (.A1(_02269_),
    .A2(_02906_),
    .B1(_02900_),
    .X(_03106_));
 sky130_fd_sc_hd__o22a_2 _08712_ (.A1(_02941_),
    .A2(_03103_),
    .B1(_03105_),
    .B2(_03106_),
    .X(\core.alu_out[23] ));
 sky130_fd_sc_hd__or4_2 _08713_ (.A(_02272_),
    .B(_02275_),
    .C(_02279_),
    .D(_02283_),
    .X(_03107_));
 sky130_fd_sc_hd__o21ai_2 _08714_ (.A1(_02278_),
    .A2(_02280_),
    .B1(_02282_),
    .Y(_03108_));
 sky130_fd_sc_hd__nor2_2 _08715_ (.A(_02273_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__or3_2 _08716_ (.A(_02271_),
    .B(_02274_),
    .C(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__o21ba_2 _08717_ (.A1(_03075_),
    .A2(_03107_),
    .B1_N(_02269_),
    .X(_03111_));
 sky130_fd_sc_hd__o211a_2 _08718_ (.A1(_03077_),
    .A2(_03107_),
    .B1(_03110_),
    .C1(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__mux2_2 _08719_ (.A0(_02412_),
    .A1(_03112_),
    .S(_02921_),
    .X(_03113_));
 sky130_fd_sc_hd__xor2_2 _08720_ (.A(_02259_),
    .B(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_2 _08721_ (.A0(_02897_),
    .A1(_02896_),
    .S(_02258_),
    .X(_03115_));
 sky130_fd_sc_hd__o21ba_2 _08722_ (.A1(_02937_),
    .A2(_03115_),
    .B1_N(_02257_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_2 _08723_ (.A0(_03114_),
    .A1(_03116_),
    .S(_02979_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_1 _08724_ (.A(_03117_),
    .X(\core.alu_out[24] ));
 sky130_fd_sc_hd__a21oi_2 _08725_ (.A1(_02254_),
    .A2(_02924_),
    .B1(_02901_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_2 _08726_ (.A(_02253_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__a31o_2 _08727_ (.A1(\core.pcpi_rs2[25] ),
    .A2(_02814_),
    .A3(_02905_),
    .B1(_02899_),
    .X(_03120_));
 sky130_fd_sc_hd__a21o_2 _08728_ (.A1(_02259_),
    .A2(_02412_),
    .B1(_02419_),
    .X(_03121_));
 sky130_fd_sc_hd__o21a_2 _08729_ (.A1(_02257_),
    .A2(_03112_),
    .B1(_02258_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_2 _08730_ (.A0(_03121_),
    .A1(_03122_),
    .S(_02912_),
    .X(_03123_));
 sky130_fd_sc_hd__xor2_2 _08731_ (.A(_02255_),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__o22a_2 _08732_ (.A1(_03119_),
    .A2(_03120_),
    .B1(_03124_),
    .B2(_02941_),
    .X(\core.alu_out[25] ));
 sky130_fd_sc_hd__a21oi_2 _08733_ (.A1(_02255_),
    .A2(_03121_),
    .B1(_02420_),
    .Y(_03125_));
 sky130_fd_sc_hd__a21oi_2 _08734_ (.A1(_02254_),
    .A2(_03122_),
    .B1(_02253_),
    .Y(_03126_));
 sky130_fd_sc_hd__mux2_2 _08735_ (.A0(_03125_),
    .A1(_03126_),
    .S(_02911_),
    .X(_03127_));
 sky130_fd_sc_hd__xor2_2 _08736_ (.A(_02266_),
    .B(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_2 _08737_ (.A0(_02902_),
    .A1(_02897_),
    .S(_02264_),
    .X(_03129_));
 sky130_fd_sc_hd__o21ba_2 _08738_ (.A1(_02937_),
    .A2(_03129_),
    .B1_N(_02265_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_2 _08739_ (.A0(_03128_),
    .A1(_03130_),
    .S(_02979_),
    .X(_03131_));
 sky130_fd_sc_hd__buf_1 _08740_ (.A(_03131_),
    .X(\core.alu_out[26] ));
 sky130_fd_sc_hd__nor2_2 _08741_ (.A(_02264_),
    .B(_03126_),
    .Y(_03132_));
 sky130_fd_sc_hd__o211ai_2 _08742_ (.A1(_02266_),
    .A2(_03125_),
    .B1(_02423_),
    .C1(_02942_),
    .Y(_03133_));
 sky130_fd_sc_hd__o31a_2 _08743_ (.A1(_02942_),
    .A2(_02265_),
    .A3(_03132_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__xnor2_2 _08744_ (.A(_02263_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_2 _08745_ (.A(\core.pcpi_rs2[27] ),
    .B(_02838_),
    .Y(_03136_));
 sky130_fd_sc_hd__a21oi_2 _08746_ (.A1(_03136_),
    .A2(_02924_),
    .B1(_02950_),
    .Y(_03137_));
 sky130_fd_sc_hd__nor2_2 _08747_ (.A(_02262_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__a21o_2 _08748_ (.A1(_02261_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_03139_));
 sky130_fd_sc_hd__o22a_2 _08749_ (.A1(_02917_),
    .A2(_03135_),
    .B1(_03138_),
    .B2(_03139_),
    .X(\core.alu_out[27] ));
 sky130_fd_sc_hd__o21ai_2 _08750_ (.A1(_02253_),
    .A2(_02258_),
    .B1(_02254_),
    .Y(_03140_));
 sky130_fd_sc_hd__nor2_2 _08751_ (.A(_02264_),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2_2 _08752_ (.A(_02263_),
    .B(_02266_),
    .Y(_03142_));
 sky130_fd_sc_hd__or4_2 _08753_ (.A(_02255_),
    .B(_02259_),
    .C(_03112_),
    .D(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__o311a_2 _08754_ (.A1(_02262_),
    .A2(_02265_),
    .A3(_03141_),
    .B1(_03143_),
    .C1(_03136_),
    .X(_03144_));
 sky130_fd_sc_hd__inv_2 _08755_ (.A(_02267_),
    .Y(_03145_));
 sky130_fd_sc_hd__a21bo_2 _08756_ (.A1(_03145_),
    .A2(_02412_),
    .B1_N(_02426_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_2 _08757_ (.A0(_03144_),
    .A1(_03146_),
    .S(_02942_),
    .X(_03147_));
 sky130_fd_sc_hd__xor2_2 _08758_ (.A(_02248_),
    .B(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__nor2_2 _08759_ (.A(_02245_),
    .B(_02907_),
    .Y(_03149_));
 sky130_fd_sc_hd__o21ba_2 _08760_ (.A1(_02950_),
    .A2(_03149_),
    .B1_N(_02247_),
    .X(_03150_));
 sky130_fd_sc_hd__a21o_2 _08761_ (.A1(_02245_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_03151_));
 sky130_fd_sc_hd__o22a_2 _08762_ (.A1(_02917_),
    .A2(_03148_),
    .B1(_03150_),
    .B2(_03151_),
    .X(\core.alu_out[28] ));
 sky130_fd_sc_hd__a21o_2 _08763_ (.A1(_02248_),
    .A2(_03146_),
    .B1(_02413_),
    .X(_03152_));
 sky130_fd_sc_hd__o21ba_2 _08764_ (.A1(_02247_),
    .A2(_03144_),
    .B1_N(_02245_),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_2 _08765_ (.A0(_03152_),
    .A1(_03153_),
    .S(_02921_),
    .X(_03154_));
 sky130_fd_sc_hd__xor2_2 _08766_ (.A(_02251_),
    .B(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__nand2_2 _08767_ (.A(\core.pcpi_rs2[29] ),
    .B(_02414_),
    .Y(_03156_));
 sky130_fd_sc_hd__a21oi_2 _08768_ (.A1(_03156_),
    .A2(_02924_),
    .B1(_02950_),
    .Y(_03157_));
 sky130_fd_sc_hd__nor2_2 _08769_ (.A(_02250_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__a21o_2 _08770_ (.A1(_02249_),
    .A2(_02906_),
    .B1(_02953_),
    .X(_03159_));
 sky130_fd_sc_hd__o22a_2 _08771_ (.A1(_02917_),
    .A2(_03155_),
    .B1(_03158_),
    .B2(_03159_),
    .X(\core.alu_out[29] ));
 sky130_fd_sc_hd__a21oi_2 _08772_ (.A1(_03156_),
    .A2(_03153_),
    .B1(_02250_),
    .Y(_03160_));
 sky130_fd_sc_hd__or2_2 _08773_ (.A(_02942_),
    .B(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__a21o_2 _08774_ (.A1(_02251_),
    .A2(_03152_),
    .B1(_02415_),
    .X(_03162_));
 sky130_fd_sc_hd__nand2_2 _08775_ (.A(_02942_),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__a21oi_2 _08776_ (.A1(_03161_),
    .A2(_03163_),
    .B1(_02244_),
    .Y(_03164_));
 sky130_fd_sc_hd__a31o_2 _08777_ (.A1(_02244_),
    .A2(_03161_),
    .A3(_03163_),
    .B1(_02917_),
    .X(_03165_));
 sky130_fd_sc_hd__o21ba_2 _08778_ (.A1(_02241_),
    .A2(_02907_),
    .B1_N(_02895_),
    .X(_03166_));
 sky130_fd_sc_hd__a2bb2o_2 _08779_ (.A1_N(_02243_),
    .A2_N(_03166_),
    .B1(_02905_),
    .B2(_02241_),
    .X(_03167_));
 sky130_fd_sc_hd__o22a_2 _08780_ (.A1(_03164_),
    .A2(_03165_),
    .B1(_03167_),
    .B2(_02900_),
    .X(\core.alu_out[30] ));
 sky130_fd_sc_hd__and2b_2 _08781_ (.A_N(_02243_),
    .B(_03160_),
    .X(_03168_));
 sky130_fd_sc_hd__a21o_2 _08782_ (.A1(_02244_),
    .A2(_03162_),
    .B1(_02417_),
    .X(_03169_));
 sky130_fd_sc_hd__nand2_2 _08783_ (.A(\core.instr_sub ),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__o31a_2 _08784_ (.A1(\core.instr_sub ),
    .A2(_02241_),
    .A3(_03168_),
    .B1(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__xnor2_2 _08785_ (.A(_02240_),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__mux2_2 _08786_ (.A0(_02898_),
    .A1(_02902_),
    .S(_02238_),
    .X(_03173_));
 sky130_fd_sc_hd__o22a_2 _08787_ (.A1(\core.pcpi_rs2[31] ),
    .A2(_02237_),
    .B1(_02937_),
    .B2(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_2 _08788_ (.A0(_03172_),
    .A1(_03174_),
    .S(_02979_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_1 _08789_ (.A(_03175_),
    .X(\core.alu_out[31] ));
 sky130_fd_sc_hd__buf_1 _08790_ (.A(_02026_),
    .X(_03176_));
 sky130_fd_sc_hd__buf_1 _08791_ (.A(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__mux2_2 _08792_ (.A0(\core.mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__buf_1 _08793_ (.A(_03178_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_2 _08794_ (.A0(\core.decoded_imm_j[15] ),
    .A1(_01358_),
    .S(_02449_),
    .X(_03179_));
 sky130_fd_sc_hd__buf_1 _08795_ (.A(_03179_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_2 _08796_ (.A0(\core.mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(_03177_),
    .X(_03180_));
 sky130_fd_sc_hd__buf_1 _08797_ (.A(_03180_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_2 _08798_ (.A0(\core.decoded_imm_j[16] ),
    .A1(_01359_),
    .S(_02449_),
    .X(_03181_));
 sky130_fd_sc_hd__buf_1 _08799_ (.A(_03181_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_2 _08800_ (.A0(\core.mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(_03177_),
    .X(_03182_));
 sky130_fd_sc_hd__buf_1 _08801_ (.A(_03182_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_2 _08802_ (.A0(\core.decoded_imm_j[17] ),
    .A1(_01360_),
    .S(_02449_),
    .X(_03183_));
 sky130_fd_sc_hd__buf_1 _08803_ (.A(_03183_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_2 _08804_ (.A0(\core.mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(_03177_),
    .X(_03184_));
 sky130_fd_sc_hd__buf_1 _08805_ (.A(_03184_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_2 _08806_ (.A0(\core.decoded_imm_j[18] ),
    .A1(_01361_),
    .S(_02449_),
    .X(_03185_));
 sky130_fd_sc_hd__buf_1 _08807_ (.A(_03185_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_2 _08808_ (.A0(\core.mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(_03177_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_1 _08809_ (.A(_03186_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_2 _08810_ (.A0(\core.decoded_imm_j[19] ),
    .A1(_01362_),
    .S(_02449_),
    .X(_03187_));
 sky130_fd_sc_hd__buf_1 _08811_ (.A(_03187_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_2 _08812_ (.A0(\core.mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(_03177_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_1 _08813_ (.A(_03188_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_2 _08814_ (.A0(\core.decoded_imm_j[11] ),
    .A1(_01363_),
    .S(_02449_),
    .X(_03189_));
 sky130_fd_sc_hd__buf_1 _08815_ (.A(_03189_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_2 _08816_ (.A0(\core.mem_rdata_q[21] ),
    .A1(mem_rdata[21]),
    .S(_03177_),
    .X(_03190_));
 sky130_fd_sc_hd__buf_1 _08817_ (.A(_03190_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_2 _08818_ (.A0(\core.decoded_imm_j[1] ),
    .A1(_01364_),
    .S(_02449_),
    .X(_03191_));
 sky130_fd_sc_hd__buf_1 _08819_ (.A(_03191_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_2 _08820_ (.A0(\core.mem_rdata_q[22] ),
    .A1(mem_rdata[22]),
    .S(_03177_),
    .X(_03192_));
 sky130_fd_sc_hd__buf_1 _08821_ (.A(_03192_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_2 _08822_ (.A0(\core.decoded_imm_j[2] ),
    .A1(_01365_),
    .S(_02449_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_1 _08823_ (.A(_03193_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_2 _08824_ (.A0(\core.mem_rdata_q[23] ),
    .A1(mem_rdata[23]),
    .S(_03176_),
    .X(_03194_));
 sky130_fd_sc_hd__buf_1 _08825_ (.A(_03194_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_2 _08826_ (.A0(\core.decoded_imm_j[3] ),
    .A1(_01366_),
    .S(_02449_),
    .X(_03195_));
 sky130_fd_sc_hd__buf_1 _08827_ (.A(_03195_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_2 _08828_ (.A0(\core.mem_rdata_q[24] ),
    .A1(mem_rdata[24]),
    .S(_03176_),
    .X(_03196_));
 sky130_fd_sc_hd__buf_1 _08829_ (.A(_03196_),
    .X(_01367_));
 sky130_fd_sc_hd__buf_1 _08830_ (.A(_02448_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_2 _08831_ (.A0(\core.decoded_imm_j[4] ),
    .A1(_01367_),
    .S(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_1 _08832_ (.A(_03198_),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_2 _08833_ (.A(\core.latched_store ),
    .B(\core.latched_branch ),
    .Y(_03199_));
 sky130_fd_sc_hd__buf_1 _08834_ (.A(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__buf_1 _08835_ (.A(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__buf_1 _08836_ (.A(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__buf_1 _08837_ (.A(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_2 _08838_ (.A0(\core.reg_out[17] ),
    .A1(\core.reg_next_pc[17] ),
    .S(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__or2_2 _08839_ (.A(\core.mem_do_prefetch ),
    .B(\core.mem_do_rinst ),
    .X(_03205_));
 sky130_fd_sc_hd__buf_1 _08840_ (.A(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__buf_1 _08841_ (.A(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__mux2_2 _08842_ (.A0(_02293_),
    .A1(_03204_),
    .S(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_2 _08843_ (.A(\core.mem_state[1] ),
    .B(\core.mem_state[0] ),
    .Y(_03209_));
 sky130_fd_sc_hd__o21ai_2 _08844_ (.A1(\core.mem_do_rdata ),
    .A2(_03206_),
    .B1(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_2 _08845_ (.A(\core.mem_do_wdata ),
    .B(_03209_),
    .Y(_03211_));
 sky130_fd_sc_hd__a21o_2 _08846_ (.A1(_03210_),
    .A2(_03211_),
    .B1(_02048_),
    .X(_03212_));
 sky130_fd_sc_hd__nor2_2 _08847_ (.A(trap),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__buf_1 _08848_ (.A(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_2 _08849_ (.A0(mem_addr[17]),
    .A1(_03208_),
    .S(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__buf_1 _08850_ (.A(_03215_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_2 _08851_ (.A0(\core.reg_out[18] ),
    .A1(\core.reg_next_pc[18] ),
    .S(_03203_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_2 _08852_ (.A0(_02298_),
    .A1(_03216_),
    .S(_03207_),
    .X(_03217_));
 sky130_fd_sc_hd__mux2_2 _08853_ (.A0(mem_addr[18]),
    .A1(_03217_),
    .S(_03214_),
    .X(_03218_));
 sky130_fd_sc_hd__buf_1 _08854_ (.A(_03218_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_2 _08855_ (.A0(\core.reg_out[19] ),
    .A1(\core.reg_next_pc[19] ),
    .S(_03203_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_2 _08856_ (.A0(_02736_),
    .A1(_03219_),
    .S(_03207_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_2 _08857_ (.A0(mem_addr[19]),
    .A1(_03220_),
    .S(_03214_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_1 _08858_ (.A(_03221_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_2 _08859_ (.A0(\core.reg_out[20] ),
    .A1(\core.reg_next_pc[20] ),
    .S(_03203_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_2 _08860_ (.A0(_02277_),
    .A1(_03222_),
    .S(_03207_),
    .X(_03223_));
 sky130_fd_sc_hd__mux2_2 _08861_ (.A0(mem_addr[20]),
    .A1(_03223_),
    .S(_03214_),
    .X(_03224_));
 sky130_fd_sc_hd__buf_1 _08862_ (.A(_03224_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_2 _08863_ (.A0(\core.reg_out[21] ),
    .A1(\core.reg_next_pc[21] ),
    .S(_03203_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_2 _08864_ (.A0(_02281_),
    .A1(_03225_),
    .S(_03207_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_2 _08865_ (.A0(mem_addr[21]),
    .A1(_03226_),
    .S(_03214_),
    .X(_03227_));
 sky130_fd_sc_hd__buf_1 _08866_ (.A(_03227_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_2 _08867_ (.A0(\core.reg_out[22] ),
    .A1(\core.reg_next_pc[22] ),
    .S(_03203_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_2 _08868_ (.A0(_02408_),
    .A1(_03228_),
    .S(_03207_),
    .X(_03229_));
 sky130_fd_sc_hd__mux2_2 _08869_ (.A0(mem_addr[22]),
    .A1(_03229_),
    .S(_03214_),
    .X(_03230_));
 sky130_fd_sc_hd__buf_1 _08870_ (.A(_03230_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_2 _08871_ (.A0(\core.reg_out[23] ),
    .A1(\core.reg_next_pc[23] ),
    .S(_03203_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_2 _08872_ (.A0(_02270_),
    .A1(_03231_),
    .S(_03207_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_2 _08873_ (.A0(mem_addr[23]),
    .A1(_03232_),
    .S(_03214_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _08874_ (.A(_03233_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_2 _08875_ (.A0(\core.reg_out[24] ),
    .A1(\core.reg_next_pc[24] ),
    .S(_03203_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_2 _08876_ (.A0(_02256_),
    .A1(_03234_),
    .S(_03207_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_1 _08877_ (.A(_03213_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_2 _08878_ (.A0(mem_addr[24]),
    .A1(_03235_),
    .S(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_1 _08879_ (.A(_03237_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_2 _08880_ (.A0(\core.reg_out[25] ),
    .A1(\core.reg_next_pc[25] ),
    .S(_03203_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_2 _08881_ (.A0(_02814_),
    .A1(_03238_),
    .S(_03207_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_2 _08882_ (.A0(mem_addr[25]),
    .A1(_03239_),
    .S(_03236_),
    .X(_03240_));
 sky130_fd_sc_hd__buf_1 _08883_ (.A(_03240_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_2 _08884_ (.A0(\core.reg_out[26] ),
    .A1(\core.reg_next_pc[26] ),
    .S(_03203_),
    .X(_03241_));
 sky130_fd_sc_hd__buf_1 _08885_ (.A(_03206_),
    .X(_03242_));
 sky130_fd_sc_hd__mux2_2 _08886_ (.A0(_02422_),
    .A1(_03241_),
    .S(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__mux2_2 _08887_ (.A0(mem_addr[26]),
    .A1(_03243_),
    .S(_03236_),
    .X(_03244_));
 sky130_fd_sc_hd__buf_1 _08888_ (.A(_03244_),
    .X(_00046_));
 sky130_fd_sc_hd__buf_1 _08889_ (.A(_03202_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_2 _08890_ (.A0(\core.reg_out[27] ),
    .A1(\core.reg_next_pc[27] ),
    .S(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_2 _08891_ (.A0(_02838_),
    .A1(_03246_),
    .S(_03242_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_2 _08892_ (.A0(mem_addr[27]),
    .A1(_03247_),
    .S(_03236_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_1 _08893_ (.A(_03248_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_2 _08894_ (.A0(\core.reg_out[28] ),
    .A1(\core.reg_next_pc[28] ),
    .S(_03245_),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_2 _08895_ (.A0(_02246_),
    .A1(_03249_),
    .S(_03242_),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_2 _08896_ (.A0(mem_addr[28]),
    .A1(_03250_),
    .S(_03236_),
    .X(_03251_));
 sky130_fd_sc_hd__buf_1 _08897_ (.A(_03251_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_2 _08898_ (.A0(\core.reg_out[29] ),
    .A1(\core.reg_next_pc[29] ),
    .S(_03245_),
    .X(_03252_));
 sky130_fd_sc_hd__mux2_2 _08899_ (.A0(_02414_),
    .A1(_03252_),
    .S(_03242_),
    .X(_03253_));
 sky130_fd_sc_hd__mux2_2 _08900_ (.A0(mem_addr[29]),
    .A1(_03253_),
    .S(_03236_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_1 _08901_ (.A(_03254_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_2 _08902_ (.A0(\core.reg_out[30] ),
    .A1(\core.reg_next_pc[30] ),
    .S(_03245_),
    .X(_03255_));
 sky130_fd_sc_hd__mux2_2 _08903_ (.A0(_02242_),
    .A1(_03255_),
    .S(_03242_),
    .X(_03256_));
 sky130_fd_sc_hd__mux2_2 _08904_ (.A0(mem_addr[30]),
    .A1(_03256_),
    .S(_03236_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_1 _08905_ (.A(_03257_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_2 _08906_ (.A0(\core.reg_out[31] ),
    .A1(\core.reg_next_pc[31] ),
    .S(_03245_),
    .X(_03258_));
 sky130_fd_sc_hd__mux2_2 _08907_ (.A0(_02237_),
    .A1(_03258_),
    .S(_03242_),
    .X(_03259_));
 sky130_fd_sc_hd__mux2_2 _08908_ (.A0(mem_addr[31]),
    .A1(_03259_),
    .S(_03236_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_1 _08909_ (.A(_03260_),
    .X(_00051_));
 sky130_fd_sc_hd__nor2_2 _08910_ (.A(\core.cpu_state[4] ),
    .B(_02041_),
    .Y(_03261_));
 sky130_fd_sc_hd__buf_1 _08911_ (.A(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__or4_2 _08912_ (.A(\core.decoded_imm_j[16] ),
    .B(\core.decoded_imm_j[17] ),
    .C(\core.decoded_imm_j[18] ),
    .D(\core.decoded_imm_j[19] ),
    .X(_03263_));
 sky130_fd_sc_hd__o21ba_2 _08913_ (.A1(\core.decoded_imm_j[15] ),
    .A2(_03263_),
    .B1_N(\core.is_lui_auipc_jal ),
    .X(_03264_));
 sky130_fd_sc_hd__buf_1 _08914_ (.A(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__buf_1 _08915_ (.A(_00009_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_1 _08916_ (.A(_00007_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _08917_ (.A(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_1 _08918_ (.A(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__buf_1 _08919_ (.A(_00005_),
    .X(_03270_));
 sky130_fd_sc_hd__buf_1 _08920_ (.A(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__buf_1 _08921_ (.A(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_1 _08922_ (.A(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_1 _08923_ (.A(_00006_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_1 _08924_ (.A(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__mux4_2 _08925_ (.A0(\core.cpuregs[8][31] ),
    .A1(\core.cpuregs[9][31] ),
    .A2(\core.cpuregs[10][31] ),
    .A3(\core.cpuregs[11][31] ),
    .S0(_03273_),
    .S1(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_1 _08926_ (.A(_00006_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_1 _08927_ (.A(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__buf_1 _08928_ (.A(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_1 _08929_ (.A(_03270_),
    .X(_03280_));
 sky130_fd_sc_hd__buf_1 _08930_ (.A(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_2 _08931_ (.A0(\core.cpuregs[14][31] ),
    .A1(\core.cpuregs[15][31] ),
    .S(_03281_),
    .X(_03282_));
 sky130_fd_sc_hd__inv_2 _08932_ (.A(_00006_),
    .Y(_03283_));
 sky130_fd_sc_hd__buf_1 _08933_ (.A(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__buf_1 _08934_ (.A(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_2 _08935_ (.A0(\core.cpuregs[12][31] ),
    .A1(\core.cpuregs[13][31] ),
    .S(_03280_),
    .X(_03286_));
 sky130_fd_sc_hd__inv_2 _08936_ (.A(_00007_),
    .Y(_03287_));
 sky130_fd_sc_hd__buf_1 _08937_ (.A(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__buf_1 _08938_ (.A(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__a21o_2 _08939_ (.A1(_03285_),
    .A2(_03286_),
    .B1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a21o_2 _08940_ (.A1(_03279_),
    .A2(_03282_),
    .B1(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__buf_1 _08941_ (.A(_00008_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_2 _08942_ (.A1(_03269_),
    .A2(_03276_),
    .B1(_03291_),
    .C1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__buf_1 _08943_ (.A(_03289_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_1 _08944_ (.A(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__buf_1 _08945_ (.A(_03271_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_1 _08946_ (.A(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__buf_1 _08947_ (.A(_00006_),
    .X(_03298_));
 sky130_fd_sc_hd__buf_1 _08948_ (.A(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__mux4_2 _08949_ (.A0(\core.cpuregs[4][31] ),
    .A1(\core.cpuregs[5][31] ),
    .A2(\core.cpuregs[6][31] ),
    .A3(\core.cpuregs[7][31] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__buf_1 _08950_ (.A(_03280_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_2 _08951_ (.A0(\core.cpuregs[2][31] ),
    .A1(\core.cpuregs[3][31] ),
    .S(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__buf_1 _08952_ (.A(_03270_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_1 _08953_ (.A(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_2 _08954_ (.A0(\core.cpuregs[0][31] ),
    .A1(\core.cpuregs[1][31] ),
    .S(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__a21o_2 _08955_ (.A1(_03285_),
    .A2(_03305_),
    .B1(_03268_),
    .X(_03306_));
 sky130_fd_sc_hd__a21o_2 _08956_ (.A1(_03279_),
    .A2(_03302_),
    .B1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__inv_2 _08957_ (.A(_00008_),
    .Y(_03308_));
 sky130_fd_sc_hd__buf_1 _08958_ (.A(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__o211a_2 _08959_ (.A1(_03295_),
    .A2(_03300_),
    .B1(_03307_),
    .C1(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__or3_2 _08960_ (.A(_03266_),
    .B(_03293_),
    .C(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__inv_2 _08961_ (.A(_00009_),
    .Y(_03312_));
 sky130_fd_sc_hd__buf_1 _08962_ (.A(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__buf_1 _08963_ (.A(_00007_),
    .X(_03314_));
 sky130_fd_sc_hd__buf_1 _08964_ (.A(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_1 _08965_ (.A(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__mux4_2 _08966_ (.A0(\core.cpuregs[16][31] ),
    .A1(\core.cpuregs[17][31] ),
    .A2(\core.cpuregs[18][31] ),
    .A3(\core.cpuregs[19][31] ),
    .S0(_03297_),
    .S1(_03275_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_2 _08967_ (.A0(\core.cpuregs[22][31] ),
    .A1(\core.cpuregs[23][31] ),
    .S(_03281_),
    .X(_03318_));
 sky130_fd_sc_hd__buf_1 _08968_ (.A(_03270_),
    .X(_03319_));
 sky130_fd_sc_hd__buf_1 _08969_ (.A(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_2 _08970_ (.A0(\core.cpuregs[20][31] ),
    .A1(\core.cpuregs[21][31] ),
    .S(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__a21o_2 _08971_ (.A1(_03285_),
    .A2(_03321_),
    .B1(_03289_),
    .X(_03322_));
 sky130_fd_sc_hd__a21o_2 _08972_ (.A1(_03279_),
    .A2(_03318_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__o211a_2 _08973_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03323_),
    .C1(_03309_),
    .X(_03324_));
 sky130_fd_sc_hd__mux4_2 _08974_ (.A0(\core.cpuregs[24][31] ),
    .A1(\core.cpuregs[25][31] ),
    .A2(\core.cpuregs[26][31] ),
    .A3(\core.cpuregs[27][31] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_03325_));
 sky130_fd_sc_hd__buf_1 _08975_ (.A(_03277_),
    .X(_03326_));
 sky130_fd_sc_hd__buf_1 _08976_ (.A(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_2 _08977_ (.A0(\core.cpuregs[30][31] ),
    .A1(\core.cpuregs[31][31] ),
    .S(_03301_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_1 _08978_ (.A(_03303_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_2 _08979_ (.A0(\core.cpuregs[28][31] ),
    .A1(\core.cpuregs[29][31] ),
    .S(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__buf_1 _08980_ (.A(_03287_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _08981_ (.A(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__a21o_2 _08982_ (.A1(_03285_),
    .A2(_03330_),
    .B1(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__a21o_2 _08983_ (.A1(_03327_),
    .A2(_03328_),
    .B1(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__buf_1 _08984_ (.A(_00008_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_1 _08985_ (.A(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__o211a_2 _08986_ (.A1(_03316_),
    .A2(_03325_),
    .B1(_03334_),
    .C1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__or3_2 _08987_ (.A(_03313_),
    .B(_03324_),
    .C(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__and2b_2 _08988_ (.A_N(\core.instr_lui ),
    .B(\core.is_lui_auipc_jal ),
    .X(_03339_));
 sky130_fd_sc_hd__buf_1 _08989_ (.A(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__a32o_2 _08990_ (.A1(_03265_),
    .A2(_03311_),
    .A3(_03338_),
    .B1(_03340_),
    .B2(\core.reg_pc[31] ),
    .X(_03341_));
 sky130_fd_sc_hd__nor3_2 _08991_ (.A(\core.instr_srl ),
    .B(\core.instr_srli ),
    .C(_02059_),
    .Y(_03342_));
 sky130_fd_sc_hd__buf_1 _08992_ (.A(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__buf_1 _08993_ (.A(_02099_),
    .X(_03344_));
 sky130_fd_sc_hd__o21a_2 _08994_ (.A1(_02242_),
    .A2(_03344_),
    .B1(\core.cpu_state[4] ),
    .X(_03345_));
 sky130_fd_sc_hd__o211a_2 _08995_ (.A1(_02838_),
    .A2(_02179_),
    .B1(_03343_),
    .C1(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__nand2_2 _08996_ (.A(_02242_),
    .B(\core.decoded_imm[30] ),
    .Y(_03347_));
 sky130_fd_sc_hd__and2_2 _08997_ (.A(_02414_),
    .B(\core.decoded_imm[29] ),
    .X(_03348_));
 sky130_fd_sc_hd__nor2_2 _08998_ (.A(_02414_),
    .B(\core.decoded_imm[29] ),
    .Y(_03349_));
 sky130_fd_sc_hd__nor2_2 _08999_ (.A(_02246_),
    .B(\core.decoded_imm[28] ),
    .Y(_03350_));
 sky130_fd_sc_hd__nor2_2 _09000_ (.A(_02838_),
    .B(\core.decoded_imm[27] ),
    .Y(_03351_));
 sky130_fd_sc_hd__xor2_2 _09001_ (.A(_02422_),
    .B(\core.decoded_imm[26] ),
    .X(_03352_));
 sky130_fd_sc_hd__or2_2 _09002_ (.A(_02814_),
    .B(\core.decoded_imm[25] ),
    .X(_03353_));
 sky130_fd_sc_hd__or2_2 _09003_ (.A(\core.pcpi_rs1[23] ),
    .B(\core.decoded_imm[23] ),
    .X(_03354_));
 sky130_fd_sc_hd__and3_2 _09004_ (.A(_02408_),
    .B(\core.decoded_imm[22] ),
    .C(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__a21oi_2 _09005_ (.A1(_02270_),
    .A2(\core.decoded_imm[23] ),
    .B1(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__xnor2_2 _09006_ (.A(\core.pcpi_rs1[22] ),
    .B(\core.decoded_imm[22] ),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_2 _09007_ (.A(\core.pcpi_rs1[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_2 _09008_ (.A(\core.pcpi_rs1[20] ),
    .B(\core.decoded_imm[20] ),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_2 _09009_ (.A(\core.pcpi_rs1[21] ),
    .B(\core.decoded_imm[21] ),
    .Y(_03360_));
 sky130_fd_sc_hd__a21o_2 _09010_ (.A1(_03358_),
    .A2(_03359_),
    .B1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__nand2_2 _09011_ (.A(\core.pcpi_rs1[23] ),
    .B(\core.decoded_imm[23] ),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_2 _09012_ (.A(_03362_),
    .B(_03354_),
    .Y(_03363_));
 sky130_fd_sc_hd__or2_2 _09013_ (.A(\core.pcpi_rs1[20] ),
    .B(\core.decoded_imm[20] ),
    .X(_03364_));
 sky130_fd_sc_hd__nand2_2 _09014_ (.A(_03359_),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__or2_2 _09015_ (.A(\core.pcpi_rs1[21] ),
    .B(\core.decoded_imm[21] ),
    .X(_03366_));
 sky130_fd_sc_hd__nand2_2 _09016_ (.A(_03358_),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__or4_2 _09017_ (.A(_03357_),
    .B(_03365_),
    .C(_03367_),
    .D(_03363_),
    .X(_03368_));
 sky130_fd_sc_hd__nor2_2 _09018_ (.A(\core.pcpi_rs1[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_2 _09019_ (.A(\core.pcpi_rs1[18] ),
    .B(\core.decoded_imm[18] ),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_2 _09020_ (.A(\core.pcpi_rs1[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_2 _09021_ (.A(\core.pcpi_rs1[16] ),
    .B(\core.decoded_imm[16] ),
    .Y(_03372_));
 sky130_fd_sc_hd__nor2_2 _09022_ (.A(\core.pcpi_rs1[17] ),
    .B(\core.decoded_imm[17] ),
    .Y(_03373_));
 sky130_fd_sc_hd__a21o_2 _09023_ (.A1(_03371_),
    .A2(_03372_),
    .B1(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__and2_2 _09024_ (.A(\core.pcpi_rs1[19] ),
    .B(\core.decoded_imm[19] ),
    .X(_03375_));
 sky130_fd_sc_hd__or2_2 _09025_ (.A(\core.pcpi_rs1[18] ),
    .B(\core.decoded_imm[18] ),
    .X(_03376_));
 sky130_fd_sc_hd__nand2_2 _09026_ (.A(_03370_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__or3_2 _09027_ (.A(_03375_),
    .B(_03369_),
    .C(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__nand2_2 _09028_ (.A(\core.pcpi_rs1[19] ),
    .B(\core.decoded_imm[19] ),
    .Y(_03379_));
 sky130_fd_sc_hd__o221a_2 _09029_ (.A1(_03369_),
    .A2(_03370_),
    .B1(_03374_),
    .B2(_03378_),
    .C1(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__o32a_2 _09030_ (.A1(_03357_),
    .A2(_03361_),
    .A3(_03363_),
    .B1(_03368_),
    .B2(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__or2_2 _09031_ (.A(\core.pcpi_rs1[14] ),
    .B(\core.decoded_imm[14] ),
    .X(_03382_));
 sky130_fd_sc_hd__nor2_2 _09032_ (.A(\core.pcpi_rs1[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_03383_));
 sky130_fd_sc_hd__nand2_2 _09033_ (.A(\core.pcpi_rs1[13] ),
    .B(\core.decoded_imm[13] ),
    .Y(_03384_));
 sky130_fd_sc_hd__or2b_2 _09034_ (.A(_03383_),
    .B_N(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__nand2_2 _09035_ (.A(\core.pcpi_rs1[12] ),
    .B(\core.decoded_imm[12] ),
    .Y(_03386_));
 sky130_fd_sc_hd__or2_2 _09036_ (.A(\core.pcpi_rs1[12] ),
    .B(\core.decoded_imm[12] ),
    .X(_03387_));
 sky130_fd_sc_hd__nand2_2 _09037_ (.A(_03386_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__or2_2 _09038_ (.A(_03385_),
    .B(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__xor2_2 _09039_ (.A(\core.pcpi_rs1[11] ),
    .B(\core.decoded_imm[11] ),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_2 _09040_ (.A(\core.pcpi_rs1[10] ),
    .B(\core.decoded_imm[10] ),
    .Y(_03391_));
 sky130_fd_sc_hd__or2_2 _09041_ (.A(\core.pcpi_rs1[10] ),
    .B(\core.decoded_imm[10] ),
    .X(_03392_));
 sky130_fd_sc_hd__nand3_2 _09042_ (.A(_03390_),
    .B(_03391_),
    .C(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_2 _09043_ (.A(_02331_),
    .B(\core.decoded_imm[9] ),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_2 _09044_ (.A(\core.pcpi_rs1[8] ),
    .B(\core.decoded_imm[8] ),
    .Y(_03395_));
 sky130_fd_sc_hd__nor2_2 _09045_ (.A(\core.pcpi_rs1[9] ),
    .B(\core.decoded_imm[9] ),
    .Y(_03396_));
 sky130_fd_sc_hd__a21o_2 _09046_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__o211a_2 _09047_ (.A1(\core.pcpi_rs1[11] ),
    .A2(\core.decoded_imm[11] ),
    .B1(\core.decoded_imm[10] ),
    .C1(\core.pcpi_rs1[10] ),
    .X(_03398_));
 sky130_fd_sc_hd__a21oi_2 _09048_ (.A1(_02336_),
    .A2(\core.decoded_imm[11] ),
    .B1(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__o21a_2 _09049_ (.A1(_03393_),
    .A2(_03397_),
    .B1(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__a21o_2 _09050_ (.A1(_03384_),
    .A2(_03386_),
    .B1(_03383_),
    .X(_03401_));
 sky130_fd_sc_hd__o21ai_2 _09051_ (.A1(_03389_),
    .A2(_03400_),
    .B1(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__a22o_2 _09052_ (.A1(_02306_),
    .A2(\core.decoded_imm[14] ),
    .B1(\core.decoded_imm[15] ),
    .B2(_02345_),
    .X(_03403_));
 sky130_fd_sc_hd__a21o_2 _09053_ (.A1(_03382_),
    .A2(_03402_),
    .B1(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__o21ai_2 _09054_ (.A1(_02345_),
    .A2(\core.decoded_imm[15] ),
    .B1(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__or2_2 _09055_ (.A(\core.pcpi_rs1[5] ),
    .B(\core.decoded_imm[5] ),
    .X(_03406_));
 sky130_fd_sc_hd__nand2_2 _09056_ (.A(_02388_),
    .B(\core.decoded_imm[5] ),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_2 _09057_ (.A(_03406_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand2_2 _09058_ (.A(\core.pcpi_rs1[4] ),
    .B(\core.decoded_imm[4] ),
    .Y(_03409_));
 sky130_fd_sc_hd__or2_2 _09059_ (.A(\core.pcpi_rs1[4] ),
    .B(\core.decoded_imm[4] ),
    .X(_03410_));
 sky130_fd_sc_hd__nand2_2 _09060_ (.A(_03409_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__nor2_2 _09061_ (.A(_02375_),
    .B(\core.decoded_imm[3] ),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_2 _09062_ (.A(_02372_),
    .B(\core.decoded_imm[2] ),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_2 _09063_ (.A(\core.pcpi_rs1[1] ),
    .B(\core.decoded_imm[1] ),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_2 _09064_ (.A(\core.pcpi_rs1[0] ),
    .B(\core.decoded_imm[0] ),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_2 _09065_ (.A(\core.pcpi_rs1[1] ),
    .B(\core.decoded_imm[1] ),
    .Y(_03416_));
 sky130_fd_sc_hd__o21a_2 _09066_ (.A1(_03414_),
    .A2(_03415_),
    .B1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__and2_2 _09067_ (.A(_02372_),
    .B(\core.decoded_imm[2] ),
    .X(_03418_));
 sky130_fd_sc_hd__o21ba_2 _09068_ (.A1(_03413_),
    .A2(_03417_),
    .B1_N(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__nand2_2 _09069_ (.A(_02375_),
    .B(\core.decoded_imm[3] ),
    .Y(_03420_));
 sky130_fd_sc_hd__o21a_2 _09070_ (.A1(_03412_),
    .A2(_03419_),
    .B1(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__nand2_2 _09071_ (.A(\core.pcpi_rs1[6] ),
    .B(\core.decoded_imm[6] ),
    .Y(_03422_));
 sky130_fd_sc_hd__or2_2 _09072_ (.A(\core.pcpi_rs1[6] ),
    .B(\core.decoded_imm[6] ),
    .X(_03423_));
 sky130_fd_sc_hd__nand2_2 _09073_ (.A(_03422_),
    .B(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__or2_2 _09074_ (.A(\core.pcpi_rs1[7] ),
    .B(\core.decoded_imm[7] ),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_2 _09075_ (.A(\core.pcpi_rs1[7] ),
    .B(\core.decoded_imm[7] ),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_2 _09076_ (.A(_03425_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__or2_2 _09077_ (.A(_03424_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__or4_2 _09078_ (.A(_03408_),
    .B(_03411_),
    .C(_03421_),
    .D(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__nand2_2 _09079_ (.A(_03426_),
    .B(_03422_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21bo_2 _09080_ (.A1(_03407_),
    .A2(_03409_),
    .B1_N(_03406_),
    .X(_03431_));
 sky130_fd_sc_hd__nor2_2 _09081_ (.A(_03424_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__o21ai_2 _09082_ (.A1(_03430_),
    .A2(_03432_),
    .B1(_03425_),
    .Y(_03433_));
 sky130_fd_sc_hd__or2b_2 _09083_ (.A(_03396_),
    .B_N(_03394_),
    .X(_03434_));
 sky130_fd_sc_hd__or2_2 _09084_ (.A(_02327_),
    .B(\core.decoded_imm[8] ),
    .X(_03435_));
 sky130_fd_sc_hd__nand2_2 _09085_ (.A(_03395_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__or3_2 _09086_ (.A(_03393_),
    .B(_03434_),
    .C(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__nand2_2 _09087_ (.A(\core.pcpi_rs1[14] ),
    .B(\core.decoded_imm[14] ),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_2 _09088_ (.A(_03382_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__xor2_2 _09089_ (.A(\core.pcpi_rs1[15] ),
    .B(\core.decoded_imm[15] ),
    .X(_03440_));
 sky130_fd_sc_hd__or3b_2 _09090_ (.A(_03389_),
    .B(_03439_),
    .C_N(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__a211o_2 _09091_ (.A1(_03429_),
    .A2(_03433_),
    .B1(_03437_),
    .C1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__or2_2 _09092_ (.A(\core.pcpi_rs1[16] ),
    .B(\core.decoded_imm[16] ),
    .X(_03443_));
 sky130_fd_sc_hd__and2_2 _09093_ (.A(_03372_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__and2b_2 _09094_ (.A_N(_03373_),
    .B(_03371_),
    .X(_03445_));
 sky130_fd_sc_hd__nand2_2 _09095_ (.A(_03444_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__a2111o_2 _09096_ (.A1(_03405_),
    .A2(_03442_),
    .B1(_03446_),
    .C1(_03378_),
    .D1(_03368_),
    .X(_03447_));
 sky130_fd_sc_hd__and3_2 _09097_ (.A(_03356_),
    .B(_03381_),
    .C(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__nand2_2 _09098_ (.A(_02256_),
    .B(\core.decoded_imm[24] ),
    .Y(_03449_));
 sky130_fd_sc_hd__or2_2 _09099_ (.A(\core.pcpi_rs1[24] ),
    .B(\core.decoded_imm[24] ),
    .X(_03450_));
 sky130_fd_sc_hd__nand2_2 _09100_ (.A(_03449_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_2 _09101_ (.A(_02814_),
    .B(\core.decoded_imm[25] ),
    .Y(_03452_));
 sky130_fd_sc_hd__o211ai_2 _09102_ (.A1(_03448_),
    .A2(_03451_),
    .B1(_03452_),
    .C1(_03449_),
    .Y(_03453_));
 sky130_fd_sc_hd__and3_2 _09103_ (.A(_03352_),
    .B(_03353_),
    .C(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__a21oi_2 _09104_ (.A1(_02422_),
    .A2(\core.decoded_imm[26] ),
    .B1(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_2 _09105_ (.A(_02838_),
    .B(\core.decoded_imm[27] ),
    .X(_03456_));
 sky130_fd_sc_hd__o21ba_2 _09106_ (.A1(_03351_),
    .A2(_03455_),
    .B1_N(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__and2_2 _09107_ (.A(_02246_),
    .B(\core.decoded_imm[28] ),
    .X(_03458_));
 sky130_fd_sc_hd__o21bai_2 _09108_ (.A1(_03350_),
    .A2(_03457_),
    .B1_N(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__and2b_2 _09109_ (.A_N(_03349_),
    .B(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__or2_2 _09110_ (.A(_02242_),
    .B(\core.decoded_imm[30] ),
    .X(_03461_));
 sky130_fd_sc_hd__o211ai_2 _09111_ (.A1(_03348_),
    .A2(_03460_),
    .B1(_03347_),
    .C1(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__xnor2_2 _09112_ (.A(_02237_),
    .B(\core.decoded_imm[31] ),
    .Y(_03463_));
 sky130_fd_sc_hd__a21oi_2 _09113_ (.A1(_03347_),
    .A2(_03462_),
    .B1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a31o_2 _09114_ (.A1(_03347_),
    .A2(_03462_),
    .A3(_03463_),
    .B1(_02121_),
    .X(_03465_));
 sky130_fd_sc_hd__nor2_2 _09115_ (.A(_03464_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__a211o_2 _09116_ (.A1(_03262_),
    .A2(_03341_),
    .B1(_03346_),
    .C1(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__or3_2 _09117_ (.A(\core.instr_srl ),
    .B(\core.instr_srli ),
    .C(_02059_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _09118_ (.A(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__o31a_2 _09119_ (.A1(\core.instr_sll ),
    .A2(\core.instr_slli ),
    .A3(_03469_),
    .B1(_02100_),
    .X(_03470_));
 sky130_fd_sc_hd__nor2_2 _09120_ (.A(\core.cpu_state[2] ),
    .B(\core.cpu_state[4] ),
    .Y(_03471_));
 sky130_fd_sc_hd__a2bb2o_2 _09121_ (.A1_N(_02125_),
    .A2_N(_03470_),
    .B1(_03471_),
    .B2(_02120_),
    .X(_03472_));
 sky130_fd_sc_hd__or4bb_2 _09122_ (.A(_02048_),
    .B(_03472_),
    .C_N(_02046_),
    .D_N(_02043_),
    .X(_03473_));
 sky130_fd_sc_hd__a21o_2 _09123_ (.A1(_02059_),
    .A2(_02102_),
    .B1(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_2 _09124_ (.A0(_03467_),
    .A1(_02237_),
    .S(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__buf_1 _09125_ (.A(_03475_),
    .X(_00052_));
 sky130_fd_sc_hd__nor2_2 _09126_ (.A(_02055_),
    .B(\core.count_cycle[0] ),
    .Y(_00053_));
 sky130_fd_sc_hd__buf_1 _09127_ (.A(_02049_),
    .X(_03476_));
 sky130_fd_sc_hd__a21oi_2 _09128_ (.A1(\core.count_cycle[0] ),
    .A2(\core.count_cycle[1] ),
    .B1(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__o21a_2 _09129_ (.A1(\core.count_cycle[0] ),
    .A2(\core.count_cycle[1] ),
    .B1(_03477_),
    .X(_00054_));
 sky130_fd_sc_hd__and3_2 _09130_ (.A(\core.count_cycle[0] ),
    .B(\core.count_cycle[1] ),
    .C(\core.count_cycle[2] ),
    .X(_03478_));
 sky130_fd_sc_hd__a21o_2 _09131_ (.A1(\core.count_cycle[0] ),
    .A2(\core.count_cycle[1] ),
    .B1(\core.count_cycle[2] ),
    .X(_03479_));
 sky130_fd_sc_hd__and3b_2 _09132_ (.A_N(_03478_),
    .B(_03479_),
    .C(_02082_),
    .X(_03480_));
 sky130_fd_sc_hd__buf_1 _09133_ (.A(_03480_),
    .X(_00055_));
 sky130_fd_sc_hd__and4_2 _09134_ (.A(\core.count_cycle[0] ),
    .B(\core.count_cycle[1] ),
    .C(\core.count_cycle[2] ),
    .D(\core.count_cycle[3] ),
    .X(_03481_));
 sky130_fd_sc_hd__buf_1 _09135_ (.A(_02052_),
    .X(_03482_));
 sky130_fd_sc_hd__o21ai_2 _09136_ (.A1(\core.count_cycle[3] ),
    .A2(_03478_),
    .B1(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__nor2_2 _09137_ (.A(_03481_),
    .B(_03483_),
    .Y(_00056_));
 sky130_fd_sc_hd__a21oi_2 _09138_ (.A1(\core.count_cycle[4] ),
    .A2(_03481_),
    .B1(_03476_),
    .Y(_03484_));
 sky130_fd_sc_hd__o21a_2 _09139_ (.A1(\core.count_cycle[4] ),
    .A2(_03481_),
    .B1(_03484_),
    .X(_00057_));
 sky130_fd_sc_hd__and3_2 _09140_ (.A(\core.count_cycle[4] ),
    .B(\core.count_cycle[5] ),
    .C(_03481_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _09141_ (.A(_02052_),
    .X(_03486_));
 sky130_fd_sc_hd__a21o_2 _09142_ (.A1(\core.count_cycle[4] ),
    .A2(_03481_),
    .B1(\core.count_cycle[5] ),
    .X(_03487_));
 sky130_fd_sc_hd__and3b_2 _09143_ (.A_N(_03485_),
    .B(_03486_),
    .C(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__buf_1 _09144_ (.A(_03488_),
    .X(_00058_));
 sky130_fd_sc_hd__and4_2 _09145_ (.A(\core.count_cycle[4] ),
    .B(\core.count_cycle[5] ),
    .C(\core.count_cycle[6] ),
    .D(_03481_),
    .X(_03489_));
 sky130_fd_sc_hd__or2_2 _09146_ (.A(\core.count_cycle[6] ),
    .B(_03485_),
    .X(_03490_));
 sky130_fd_sc_hd__and3b_2 _09147_ (.A_N(_03489_),
    .B(_03486_),
    .C(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _09148_ (.A(_03491_),
    .X(_00059_));
 sky130_fd_sc_hd__a21oi_2 _09149_ (.A1(\core.count_cycle[7] ),
    .A2(_03489_),
    .B1(_03476_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21a_2 _09150_ (.A1(\core.count_cycle[7] ),
    .A2(_03489_),
    .B1(_03492_),
    .X(_00060_));
 sky130_fd_sc_hd__and3_2 _09151_ (.A(\core.count_cycle[7] ),
    .B(\core.count_cycle[8] ),
    .C(_03489_),
    .X(_03493_));
 sky130_fd_sc_hd__a21o_2 _09152_ (.A1(\core.count_cycle[7] ),
    .A2(_03489_),
    .B1(\core.count_cycle[8] ),
    .X(_03494_));
 sky130_fd_sc_hd__and3b_2 _09153_ (.A_N(_03493_),
    .B(_03486_),
    .C(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__buf_1 _09154_ (.A(_03495_),
    .X(_00061_));
 sky130_fd_sc_hd__and2_2 _09155_ (.A(\core.count_cycle[9] ),
    .B(_03493_),
    .X(_03496_));
 sky130_fd_sc_hd__o21ai_2 _09156_ (.A1(\core.count_cycle[9] ),
    .A2(_03493_),
    .B1(_03482_),
    .Y(_03497_));
 sky130_fd_sc_hd__nor2_2 _09157_ (.A(_03496_),
    .B(_03497_),
    .Y(_00062_));
 sky130_fd_sc_hd__buf_1 _09158_ (.A(_02049_),
    .X(_03498_));
 sky130_fd_sc_hd__and3_2 _09159_ (.A(\core.count_cycle[9] ),
    .B(\core.count_cycle[10] ),
    .C(_03493_),
    .X(_03499_));
 sky130_fd_sc_hd__nor2_2 _09160_ (.A(_03498_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__o21a_2 _09161_ (.A1(\core.count_cycle[10] ),
    .A2(_03496_),
    .B1(_03500_),
    .X(_00063_));
 sky130_fd_sc_hd__a21o_2 _09162_ (.A1(\core.count_cycle[11] ),
    .A2(_03499_),
    .B1(_02054_),
    .X(_03501_));
 sky130_fd_sc_hd__o21ba_2 _09163_ (.A1(\core.count_cycle[11] ),
    .A2(_03499_),
    .B1_N(_03501_),
    .X(_00064_));
 sky130_fd_sc_hd__and3_2 _09164_ (.A(\core.count_cycle[11] ),
    .B(\core.count_cycle[12] ),
    .C(_03499_),
    .X(_03502_));
 sky130_fd_sc_hd__and2_2 _09165_ (.A(\core.count_cycle[8] ),
    .B(\core.count_cycle[9] ),
    .X(_03503_));
 sky130_fd_sc_hd__and4_2 _09166_ (.A(\core.count_cycle[7] ),
    .B(\core.count_cycle[10] ),
    .C(_03489_),
    .D(_03503_),
    .X(_03504_));
 sky130_fd_sc_hd__a21o_2 _09167_ (.A1(\core.count_cycle[11] ),
    .A2(_03504_),
    .B1(\core.count_cycle[12] ),
    .X(_03505_));
 sky130_fd_sc_hd__and3b_2 _09168_ (.A_N(_03502_),
    .B(_03486_),
    .C(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__buf_1 _09169_ (.A(_03506_),
    .X(_00065_));
 sky130_fd_sc_hd__and4_2 _09170_ (.A(\core.count_cycle[11] ),
    .B(\core.count_cycle[12] ),
    .C(\core.count_cycle[13] ),
    .D(_03504_),
    .X(_03507_));
 sky130_fd_sc_hd__or2_2 _09171_ (.A(\core.count_cycle[13] ),
    .B(_03502_),
    .X(_03508_));
 sky130_fd_sc_hd__and3b_2 _09172_ (.A_N(_03507_),
    .B(_03486_),
    .C(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__buf_1 _09173_ (.A(_03509_),
    .X(_00066_));
 sky130_fd_sc_hd__and3_2 _09174_ (.A(\core.count_cycle[13] ),
    .B(\core.count_cycle[14] ),
    .C(_03502_),
    .X(_03510_));
 sky130_fd_sc_hd__nor2_2 _09175_ (.A(_03498_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__o21a_2 _09176_ (.A1(\core.count_cycle[14] ),
    .A2(_03507_),
    .B1(_03511_),
    .X(_00067_));
 sky130_fd_sc_hd__and2_2 _09177_ (.A(\core.count_cycle[15] ),
    .B(_03510_),
    .X(_03512_));
 sky130_fd_sc_hd__or2_2 _09178_ (.A(\core.count_cycle[15] ),
    .B(_03510_),
    .X(_03513_));
 sky130_fd_sc_hd__and3b_2 _09179_ (.A_N(_03512_),
    .B(_03486_),
    .C(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__buf_1 _09180_ (.A(_03514_),
    .X(_00068_));
 sky130_fd_sc_hd__and4_2 _09181_ (.A(\core.count_cycle[14] ),
    .B(\core.count_cycle[15] ),
    .C(\core.count_cycle[16] ),
    .D(_03507_),
    .X(_03515_));
 sky130_fd_sc_hd__or2_2 _09182_ (.A(\core.count_cycle[16] ),
    .B(_03512_),
    .X(_03516_));
 sky130_fd_sc_hd__and3b_2 _09183_ (.A_N(_03515_),
    .B(_03486_),
    .C(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__buf_1 _09184_ (.A(_03517_),
    .X(_00069_));
 sky130_fd_sc_hd__and2_2 _09185_ (.A(\core.count_cycle[17] ),
    .B(_03515_),
    .X(_03518_));
 sky130_fd_sc_hd__or2_2 _09186_ (.A(\core.count_cycle[17] ),
    .B(_03515_),
    .X(_03519_));
 sky130_fd_sc_hd__and3b_2 _09187_ (.A_N(_03518_),
    .B(_03486_),
    .C(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__buf_1 _09188_ (.A(_03520_),
    .X(_00070_));
 sky130_fd_sc_hd__nor2_2 _09189_ (.A(\core.count_cycle[18] ),
    .B(_03518_),
    .Y(_03521_));
 sky130_fd_sc_hd__and3_2 _09190_ (.A(\core.count_cycle[17] ),
    .B(\core.count_cycle[18] ),
    .C(_03515_),
    .X(_03522_));
 sky130_fd_sc_hd__nor3_2 _09191_ (.A(_03476_),
    .B(_03521_),
    .C(_03522_),
    .Y(_00071_));
 sky130_fd_sc_hd__and4_2 _09192_ (.A(\core.count_cycle[17] ),
    .B(\core.count_cycle[18] ),
    .C(\core.count_cycle[19] ),
    .D(_03515_),
    .X(_03523_));
 sky130_fd_sc_hd__buf_1 _09193_ (.A(_02052_),
    .X(_03524_));
 sky130_fd_sc_hd__or2_2 _09194_ (.A(\core.count_cycle[19] ),
    .B(_03522_),
    .X(_03525_));
 sky130_fd_sc_hd__and3b_2 _09195_ (.A_N(_03523_),
    .B(_03524_),
    .C(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__buf_1 _09196_ (.A(_03526_),
    .X(_00072_));
 sky130_fd_sc_hd__and4_2 _09197_ (.A(\core.count_cycle[16] ),
    .B(\core.count_cycle[17] ),
    .C(\core.count_cycle[18] ),
    .D(_03512_),
    .X(_03527_));
 sky130_fd_sc_hd__a31o_2 _09198_ (.A1(\core.count_cycle[19] ),
    .A2(\core.count_cycle[20] ),
    .A3(_03527_),
    .B1(_02054_),
    .X(_03528_));
 sky130_fd_sc_hd__o21ba_2 _09199_ (.A1(\core.count_cycle[20] ),
    .A2(_03523_),
    .B1_N(_03528_),
    .X(_00073_));
 sky130_fd_sc_hd__and4_2 _09200_ (.A(\core.count_cycle[19] ),
    .B(\core.count_cycle[20] ),
    .C(\core.count_cycle[21] ),
    .D(_03527_),
    .X(_03529_));
 sky130_fd_sc_hd__a21o_2 _09201_ (.A1(\core.count_cycle[20] ),
    .A2(_03523_),
    .B1(\core.count_cycle[21] ),
    .X(_03530_));
 sky130_fd_sc_hd__and3b_2 _09202_ (.A_N(_03529_),
    .B(_03530_),
    .C(_02082_),
    .X(_03531_));
 sky130_fd_sc_hd__buf_1 _09203_ (.A(_03531_),
    .X(_00074_));
 sky130_fd_sc_hd__and2_2 _09204_ (.A(\core.count_cycle[21] ),
    .B(\core.count_cycle[22] ),
    .X(_03532_));
 sky130_fd_sc_hd__a31o_2 _09205_ (.A1(\core.count_cycle[20] ),
    .A2(_03523_),
    .A3(_03532_),
    .B1(_02049_),
    .X(_03533_));
 sky130_fd_sc_hd__o21ba_2 _09206_ (.A1(\core.count_cycle[22] ),
    .A2(_03529_),
    .B1_N(_03533_),
    .X(_00075_));
 sky130_fd_sc_hd__and4_2 _09207_ (.A(\core.count_cycle[20] ),
    .B(\core.count_cycle[23] ),
    .C(_03523_),
    .D(_03532_),
    .X(_03534_));
 sky130_fd_sc_hd__a31o_2 _09208_ (.A1(\core.count_cycle[20] ),
    .A2(_03523_),
    .A3(_03532_),
    .B1(\core.count_cycle[23] ),
    .X(_03535_));
 sky130_fd_sc_hd__and3b_2 _09209_ (.A_N(_03534_),
    .B(_03524_),
    .C(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__buf_1 _09210_ (.A(_03536_),
    .X(_00076_));
 sky130_fd_sc_hd__and4_2 _09211_ (.A(\core.count_cycle[22] ),
    .B(\core.count_cycle[23] ),
    .C(\core.count_cycle[24] ),
    .D(_03529_),
    .X(_03537_));
 sky130_fd_sc_hd__nor2_2 _09212_ (.A(_03498_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__o21a_2 _09213_ (.A1(\core.count_cycle[24] ),
    .A2(_03534_),
    .B1(_03538_),
    .X(_00077_));
 sky130_fd_sc_hd__and2_2 _09214_ (.A(\core.count_cycle[24] ),
    .B(\core.count_cycle[25] ),
    .X(_03539_));
 sky130_fd_sc_hd__a21oi_2 _09215_ (.A1(_03534_),
    .A2(_03539_),
    .B1(_03498_),
    .Y(_03540_));
 sky130_fd_sc_hd__o21a_2 _09216_ (.A1(\core.count_cycle[25] ),
    .A2(_03537_),
    .B1(_03540_),
    .X(_00078_));
 sky130_fd_sc_hd__and3_2 _09217_ (.A(\core.count_cycle[25] ),
    .B(\core.count_cycle[26] ),
    .C(_03537_),
    .X(_03541_));
 sky130_fd_sc_hd__a21o_2 _09218_ (.A1(_03534_),
    .A2(_03539_),
    .B1(\core.count_cycle[26] ),
    .X(_03542_));
 sky130_fd_sc_hd__and3b_2 _09219_ (.A_N(_03541_),
    .B(_03524_),
    .C(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__buf_1 _09220_ (.A(_03543_),
    .X(_00079_));
 sky130_fd_sc_hd__and4_2 _09221_ (.A(\core.count_cycle[25] ),
    .B(\core.count_cycle[26] ),
    .C(\core.count_cycle[27] ),
    .D(_03537_),
    .X(_03544_));
 sky130_fd_sc_hd__nor2_2 _09222_ (.A(_03498_),
    .B(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__o21a_2 _09223_ (.A1(\core.count_cycle[27] ),
    .A2(_03541_),
    .B1(_03545_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_1 _09224_ (.A(_02052_),
    .X(_03546_));
 sky130_fd_sc_hd__and4_2 _09225_ (.A(\core.count_cycle[26] ),
    .B(\core.count_cycle[27] ),
    .C(_03534_),
    .D(_03539_),
    .X(_03547_));
 sky130_fd_sc_hd__or2_2 _09226_ (.A(\core.count_cycle[28] ),
    .B(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__nand2_2 _09227_ (.A(\core.count_cycle[28] ),
    .B(_03544_),
    .Y(_03549_));
 sky130_fd_sc_hd__and3_2 _09228_ (.A(_03546_),
    .B(_03548_),
    .C(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_1 _09229_ (.A(_03550_),
    .X(_00081_));
 sky130_fd_sc_hd__inv_2 _09230_ (.A(\core.count_cycle[29] ),
    .Y(_03551_));
 sky130_fd_sc_hd__and2_2 _09231_ (.A(\core.count_cycle[28] ),
    .B(\core.count_cycle[29] ),
    .X(_03552_));
 sky130_fd_sc_hd__and2_2 _09232_ (.A(_03544_),
    .B(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a211oi_2 _09233_ (.A1(_03551_),
    .A2(_03549_),
    .B1(_03553_),
    .C1(_03476_),
    .Y(_00082_));
 sky130_fd_sc_hd__and3_2 _09234_ (.A(\core.count_cycle[30] ),
    .B(_03544_),
    .C(_03552_),
    .X(_03554_));
 sky130_fd_sc_hd__or2_2 _09235_ (.A(\core.count_cycle[30] ),
    .B(_03553_),
    .X(_03555_));
 sky130_fd_sc_hd__and3b_2 _09236_ (.A_N(_03554_),
    .B(_03524_),
    .C(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_1 _09237_ (.A(_03556_),
    .X(_00083_));
 sky130_fd_sc_hd__buf_1 _09238_ (.A(_02049_),
    .X(_03557_));
 sky130_fd_sc_hd__and4_2 _09239_ (.A(\core.count_cycle[30] ),
    .B(\core.count_cycle[31] ),
    .C(_03544_),
    .D(_03552_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_2 _09240_ (.A(_03557_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__o21a_2 _09241_ (.A1(\core.count_cycle[31] ),
    .A2(_03554_),
    .B1(_03559_),
    .X(_00084_));
 sky130_fd_sc_hd__and4_2 _09242_ (.A(\core.count_cycle[30] ),
    .B(\core.count_cycle[31] ),
    .C(_03547_),
    .D(_03552_),
    .X(_03560_));
 sky130_fd_sc_hd__or2_2 _09243_ (.A(\core.count_cycle[32] ),
    .B(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_2 _09244_ (.A(\core.count_cycle[32] ),
    .B(_03558_),
    .Y(_03562_));
 sky130_fd_sc_hd__and3_2 _09245_ (.A(_03546_),
    .B(_03561_),
    .C(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__buf_1 _09246_ (.A(_03563_),
    .X(_00085_));
 sky130_fd_sc_hd__inv_2 _09247_ (.A(\core.count_cycle[33] ),
    .Y(_03564_));
 sky130_fd_sc_hd__and2_2 _09248_ (.A(\core.count_cycle[32] ),
    .B(\core.count_cycle[33] ),
    .X(_03565_));
 sky130_fd_sc_hd__and2_2 _09249_ (.A(_03558_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__a211oi_2 _09250_ (.A1(_03564_),
    .A2(_03562_),
    .B1(_03566_),
    .C1(_03476_),
    .Y(_00086_));
 sky130_fd_sc_hd__and3_2 _09251_ (.A(\core.count_cycle[34] ),
    .B(_03558_),
    .C(_03565_),
    .X(_03567_));
 sky130_fd_sc_hd__nor2_2 _09252_ (.A(_03557_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__o21a_2 _09253_ (.A1(\core.count_cycle[34] ),
    .A2(_03566_),
    .B1(_03568_),
    .X(_00087_));
 sky130_fd_sc_hd__and4_2 _09254_ (.A(\core.count_cycle[34] ),
    .B(\core.count_cycle[35] ),
    .C(_03558_),
    .D(_03565_),
    .X(_03569_));
 sky130_fd_sc_hd__nor2_2 _09255_ (.A(_03557_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__o21a_2 _09256_ (.A1(\core.count_cycle[35] ),
    .A2(_03567_),
    .B1(_03570_),
    .X(_00088_));
 sky130_fd_sc_hd__buf_1 _09257_ (.A(_02052_),
    .X(_03571_));
 sky130_fd_sc_hd__and4_2 _09258_ (.A(\core.count_cycle[34] ),
    .B(\core.count_cycle[35] ),
    .C(_03560_),
    .D(_03565_),
    .X(_03572_));
 sky130_fd_sc_hd__or2_2 _09259_ (.A(\core.count_cycle[36] ),
    .B(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__nand2_2 _09260_ (.A(\core.count_cycle[36] ),
    .B(_03569_),
    .Y(_03574_));
 sky130_fd_sc_hd__and3_2 _09261_ (.A(_03571_),
    .B(_03573_),
    .C(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__buf_1 _09262_ (.A(_03575_),
    .X(_00089_));
 sky130_fd_sc_hd__inv_2 _09263_ (.A(\core.count_cycle[37] ),
    .Y(_03576_));
 sky130_fd_sc_hd__and2_2 _09264_ (.A(\core.count_cycle[36] ),
    .B(\core.count_cycle[37] ),
    .X(_03577_));
 sky130_fd_sc_hd__and2_2 _09265_ (.A(_03569_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__a211oi_2 _09266_ (.A1(_03576_),
    .A2(_03574_),
    .B1(_03578_),
    .C1(_03476_),
    .Y(_00090_));
 sky130_fd_sc_hd__and3_2 _09267_ (.A(\core.count_cycle[38] ),
    .B(_03569_),
    .C(_03577_),
    .X(_03579_));
 sky130_fd_sc_hd__nor2_2 _09268_ (.A(_03557_),
    .B(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__o21a_2 _09269_ (.A1(\core.count_cycle[38] ),
    .A2(_03578_),
    .B1(_03580_),
    .X(_00091_));
 sky130_fd_sc_hd__and2_2 _09270_ (.A(\core.count_cycle[39] ),
    .B(_03579_),
    .X(_03581_));
 sky130_fd_sc_hd__buf_1 _09271_ (.A(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__nor2_2 _09272_ (.A(_03557_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__o21a_2 _09273_ (.A1(\core.count_cycle[39] ),
    .A2(_03579_),
    .B1(_03583_),
    .X(_00092_));
 sky130_fd_sc_hd__a21oi_2 _09274_ (.A1(\core.count_cycle[40] ),
    .A2(_03582_),
    .B1(_03498_),
    .Y(_03584_));
 sky130_fd_sc_hd__o21a_2 _09275_ (.A1(\core.count_cycle[40] ),
    .A2(_03582_),
    .B1(_03584_),
    .X(_00093_));
 sky130_fd_sc_hd__and4_2 _09276_ (.A(\core.count_cycle[38] ),
    .B(\core.count_cycle[39] ),
    .C(_03572_),
    .D(_03577_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_2 _09277_ (.A1(\core.count_cycle[40] ),
    .A2(_03585_),
    .B1(\core.count_cycle[41] ),
    .X(_03586_));
 sky130_fd_sc_hd__and2_2 _09278_ (.A(\core.count_cycle[40] ),
    .B(\core.count_cycle[41] ),
    .X(_03587_));
 sky130_fd_sc_hd__nand2_2 _09279_ (.A(_03582_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__and3_2 _09280_ (.A(_03571_),
    .B(_03586_),
    .C(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__buf_1 _09281_ (.A(_03589_),
    .X(_00094_));
 sky130_fd_sc_hd__inv_2 _09282_ (.A(\core.count_cycle[42] ),
    .Y(_03590_));
 sky130_fd_sc_hd__a31o_2 _09283_ (.A1(\core.count_cycle[42] ),
    .A2(_03582_),
    .A3(_03587_),
    .B1(_02049_),
    .X(_03591_));
 sky130_fd_sc_hd__a21oi_2 _09284_ (.A1(_03590_),
    .A2(_03588_),
    .B1(_03591_),
    .Y(_00095_));
 sky130_fd_sc_hd__and4_2 _09285_ (.A(\core.count_cycle[42] ),
    .B(\core.count_cycle[43] ),
    .C(_03585_),
    .D(_03587_),
    .X(_03592_));
 sky130_fd_sc_hd__a31o_2 _09286_ (.A1(\core.count_cycle[42] ),
    .A2(_03585_),
    .A3(_03587_),
    .B1(\core.count_cycle[43] ),
    .X(_03593_));
 sky130_fd_sc_hd__and3b_2 _09287_ (.A_N(_03592_),
    .B(_03524_),
    .C(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_1 _09288_ (.A(_03594_),
    .X(_00096_));
 sky130_fd_sc_hd__or2_2 _09289_ (.A(\core.count_cycle[44] ),
    .B(_03592_),
    .X(_03595_));
 sky130_fd_sc_hd__and4_2 _09290_ (.A(\core.count_cycle[42] ),
    .B(\core.count_cycle[43] ),
    .C(_03582_),
    .D(_03587_),
    .X(_03596_));
 sky130_fd_sc_hd__nand2_2 _09291_ (.A(\core.count_cycle[44] ),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__and3_2 _09292_ (.A(_03571_),
    .B(_03595_),
    .C(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__buf_1 _09293_ (.A(_03598_),
    .X(_00097_));
 sky130_fd_sc_hd__inv_2 _09294_ (.A(\core.count_cycle[45] ),
    .Y(_03599_));
 sky130_fd_sc_hd__and2_2 _09295_ (.A(\core.count_cycle[44] ),
    .B(\core.count_cycle[45] ),
    .X(_03600_));
 sky130_fd_sc_hd__a221oi_2 _09296_ (.A1(_03599_),
    .A2(_03597_),
    .B1(_03600_),
    .B2(_03596_),
    .C1(_03476_),
    .Y(_00098_));
 sky130_fd_sc_hd__and3_2 _09297_ (.A(\core.count_cycle[46] ),
    .B(_03592_),
    .C(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__a21o_2 _09298_ (.A1(_03592_),
    .A2(_03600_),
    .B1(\core.count_cycle[46] ),
    .X(_03602_));
 sky130_fd_sc_hd__and3b_2 _09299_ (.A_N(_03601_),
    .B(_03524_),
    .C(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__buf_1 _09300_ (.A(_03603_),
    .X(_00099_));
 sky130_fd_sc_hd__and4_2 _09301_ (.A(\core.count_cycle[46] ),
    .B(\core.count_cycle[47] ),
    .C(_03592_),
    .D(_03600_),
    .X(_03604_));
 sky130_fd_sc_hd__or2_2 _09302_ (.A(\core.count_cycle[47] ),
    .B(_03601_),
    .X(_03605_));
 sky130_fd_sc_hd__and3b_2 _09303_ (.A_N(_03604_),
    .B(_03524_),
    .C(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__buf_1 _09304_ (.A(_03606_),
    .X(_00100_));
 sky130_fd_sc_hd__or2_2 _09305_ (.A(\core.count_cycle[48] ),
    .B(_03604_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_2 _09306_ (.A(\core.count_cycle[48] ),
    .B(_03604_),
    .Y(_03608_));
 sky130_fd_sc_hd__and3_2 _09307_ (.A(_03571_),
    .B(_03607_),
    .C(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__buf_1 _09308_ (.A(_03609_),
    .X(_00101_));
 sky130_fd_sc_hd__and2_2 _09309_ (.A(\core.count_cycle[48] ),
    .B(\core.count_cycle[49] ),
    .X(_03610_));
 sky130_fd_sc_hd__and2_2 _09310_ (.A(_03604_),
    .B(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__a21o_2 _09311_ (.A1(\core.count_cycle[48] ),
    .A2(_03604_),
    .B1(\core.count_cycle[49] ),
    .X(_03612_));
 sky130_fd_sc_hd__and3b_2 _09312_ (.A_N(_03611_),
    .B(_03524_),
    .C(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__buf_1 _09313_ (.A(_03613_),
    .X(_00102_));
 sky130_fd_sc_hd__and3_2 _09314_ (.A(\core.count_cycle[50] ),
    .B(_03604_),
    .C(_03610_),
    .X(_03614_));
 sky130_fd_sc_hd__or2_2 _09315_ (.A(\core.count_cycle[50] ),
    .B(_03611_),
    .X(_03615_));
 sky130_fd_sc_hd__and3b_2 _09316_ (.A_N(_03614_),
    .B(_03524_),
    .C(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__buf_1 _09317_ (.A(_03616_),
    .X(_00103_));
 sky130_fd_sc_hd__and4_2 _09318_ (.A(\core.count_cycle[50] ),
    .B(\core.count_cycle[51] ),
    .C(_03604_),
    .D(_03610_),
    .X(_03617_));
 sky130_fd_sc_hd__or2_2 _09319_ (.A(\core.count_cycle[51] ),
    .B(_03614_),
    .X(_03618_));
 sky130_fd_sc_hd__and3b_2 _09320_ (.A_N(_03617_),
    .B(_03524_),
    .C(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__buf_1 _09321_ (.A(_03619_),
    .X(_00104_));
 sky130_fd_sc_hd__and2_2 _09322_ (.A(\core.count_cycle[52] ),
    .B(_03617_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _09323_ (.A(_02024_),
    .X(_03621_));
 sky130_fd_sc_hd__or2_2 _09324_ (.A(\core.count_cycle[52] ),
    .B(_03617_),
    .X(_03622_));
 sky130_fd_sc_hd__and3b_2 _09325_ (.A_N(_03620_),
    .B(_03621_),
    .C(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__buf_1 _09326_ (.A(_03623_),
    .X(_00105_));
 sky130_fd_sc_hd__or2_2 _09327_ (.A(\core.count_cycle[53] ),
    .B(_03620_),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_2 _09328_ (.A(\core.count_cycle[53] ),
    .B(_03620_),
    .Y(_03625_));
 sky130_fd_sc_hd__and3_2 _09329_ (.A(_03571_),
    .B(_03624_),
    .C(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_1 _09330_ (.A(_03626_),
    .X(_00106_));
 sky130_fd_sc_hd__inv_2 _09331_ (.A(\core.count_cycle[54] ),
    .Y(_03627_));
 sky130_fd_sc_hd__and2_2 _09332_ (.A(\core.count_cycle[53] ),
    .B(\core.count_cycle[54] ),
    .X(_03628_));
 sky130_fd_sc_hd__and3_2 _09333_ (.A(\core.count_cycle[52] ),
    .B(_03617_),
    .C(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__a211oi_2 _09334_ (.A1(_03627_),
    .A2(_03625_),
    .B1(_03629_),
    .C1(_03476_),
    .Y(_00107_));
 sky130_fd_sc_hd__and2_2 _09335_ (.A(\core.count_cycle[55] ),
    .B(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__or2_2 _09336_ (.A(\core.count_cycle[55] ),
    .B(_03629_),
    .X(_03631_));
 sky130_fd_sc_hd__and3b_2 _09337_ (.A_N(_03630_),
    .B(_03621_),
    .C(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__buf_1 _09338_ (.A(_03632_),
    .X(_00108_));
 sky130_fd_sc_hd__and3_2 _09339_ (.A(\core.count_cycle[55] ),
    .B(\core.count_cycle[56] ),
    .C(_03629_),
    .X(_03633_));
 sky130_fd_sc_hd__or2_2 _09340_ (.A(\core.count_cycle[56] ),
    .B(_03630_),
    .X(_03634_));
 sky130_fd_sc_hd__and3b_2 _09341_ (.A_N(_03633_),
    .B(_03621_),
    .C(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _09342_ (.A(_03635_),
    .X(_00109_));
 sky130_fd_sc_hd__or2_2 _09343_ (.A(\core.count_cycle[57] ),
    .B(_03633_),
    .X(_03636_));
 sky130_fd_sc_hd__nand2_2 _09344_ (.A(\core.count_cycle[57] ),
    .B(_03633_),
    .Y(_03637_));
 sky130_fd_sc_hd__and3_2 _09345_ (.A(_03571_),
    .B(_03636_),
    .C(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_1 _09346_ (.A(_03638_),
    .X(_00110_));
 sky130_fd_sc_hd__inv_2 _09347_ (.A(\core.count_cycle[58] ),
    .Y(_03639_));
 sky130_fd_sc_hd__and4_2 _09348_ (.A(\core.count_cycle[55] ),
    .B(\core.count_cycle[56] ),
    .C(\core.count_cycle[57] ),
    .D(\core.count_cycle[58] ),
    .X(_03640_));
 sky130_fd_sc_hd__and4_2 _09349_ (.A(\core.count_cycle[52] ),
    .B(_03617_),
    .C(_03628_),
    .D(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__a211oi_2 _09350_ (.A1(_03639_),
    .A2(_03637_),
    .B1(_03641_),
    .C1(_03476_),
    .Y(_00111_));
 sky130_fd_sc_hd__and2_2 _09351_ (.A(\core.count_cycle[59] ),
    .B(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__or2_2 _09352_ (.A(\core.count_cycle[59] ),
    .B(_03641_),
    .X(_03643_));
 sky130_fd_sc_hd__and3b_2 _09353_ (.A_N(_03642_),
    .B(_03621_),
    .C(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_1 _09354_ (.A(_03644_),
    .X(_00112_));
 sky130_fd_sc_hd__and3_2 _09355_ (.A(\core.count_cycle[59] ),
    .B(\core.count_cycle[60] ),
    .C(_03641_),
    .X(_03645_));
 sky130_fd_sc_hd__or2_2 _09356_ (.A(\core.count_cycle[60] ),
    .B(_03642_),
    .X(_03646_));
 sky130_fd_sc_hd__and3b_2 _09357_ (.A_N(_03645_),
    .B(_03621_),
    .C(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_1 _09358_ (.A(_03647_),
    .X(_00113_));
 sky130_fd_sc_hd__or2_2 _09359_ (.A(\core.count_cycle[61] ),
    .B(_03645_),
    .X(_03648_));
 sky130_fd_sc_hd__nand2_2 _09360_ (.A(\core.count_cycle[61] ),
    .B(_03645_),
    .Y(_03649_));
 sky130_fd_sc_hd__and3_2 _09361_ (.A(_03571_),
    .B(_03648_),
    .C(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__buf_1 _09362_ (.A(_03650_),
    .X(_00114_));
 sky130_fd_sc_hd__a21o_2 _09363_ (.A1(\core.count_cycle[61] ),
    .A2(_03645_),
    .B1(\core.count_cycle[62] ),
    .X(_03651_));
 sky130_fd_sc_hd__nand3_2 _09364_ (.A(\core.count_cycle[61] ),
    .B(\core.count_cycle[62] ),
    .C(_03645_),
    .Y(_03652_));
 sky130_fd_sc_hd__and3_2 _09365_ (.A(_03571_),
    .B(_03651_),
    .C(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__buf_1 _09366_ (.A(_03653_),
    .X(_00115_));
 sky130_fd_sc_hd__xor2_2 _09367_ (.A(\core.count_cycle[63] ),
    .B(_03652_),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_2 _09368_ (.A(_02055_),
    .B(_03654_),
    .Y(_00116_));
 sky130_fd_sc_hd__buf_1 _09369_ (.A(_02079_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_1 _09370_ (.A(\core.latched_stalu ),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_2 _09371_ (.A0(\core.reg_out[1] ),
    .A1(\core.alu_out_q[1] ),
    .S(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_2 _09372_ (.A0(_03657_),
    .A1(\core.reg_next_pc[1] ),
    .S(_03200_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _09373_ (.A(\core.decoder_trigger ),
    .X(_03659_));
 sky130_fd_sc_hd__and2_2 _09374_ (.A(\core.instr_jal ),
    .B(\core.decoded_imm_j[1] ),
    .X(_03660_));
 sky130_fd_sc_hd__nand2_2 _09375_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__nor2_2 _09376_ (.A(_03658_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__buf_1 _09377_ (.A(_02110_),
    .X(_03663_));
 sky130_fd_sc_hd__a21o_2 _09378_ (.A1(_03658_),
    .A2(_03661_),
    .B1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__buf_1 _09379_ (.A(_03486_),
    .X(_03665_));
 sky130_fd_sc_hd__o221a_2 _09380_ (.A1(_03655_),
    .A2(\core.reg_next_pc[1] ),
    .B1(_03662_),
    .B2(_03664_),
    .C1(_03665_),
    .X(_00117_));
 sky130_fd_sc_hd__inv_2 _09381_ (.A(\core.instr_jal ),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_2 _09382_ (.A(\core.decoder_trigger ),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__mux2_2 _09383_ (.A0(\core.reg_out[2] ),
    .A1(\core.alu_out_q[2] ),
    .S(\core.latched_stalu ),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_2 _09384_ (.A0(_03668_),
    .A1(\core.reg_next_pc[2] ),
    .S(_03199_),
    .X(_03669_));
 sky130_fd_sc_hd__buf_1 _09385_ (.A(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o21ai_2 _09386_ (.A1(_03667_),
    .A2(_03670_),
    .B1(_02080_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_2 _09387_ (.A(\core.decoder_trigger ),
    .B(\core.instr_jal ),
    .Y(_03672_));
 sky130_fd_sc_hd__inv_2 _09388_ (.A(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__xor2_2 _09389_ (.A(\core.decoded_imm_j[2] ),
    .B(_03670_),
    .X(_03674_));
 sky130_fd_sc_hd__a21o_2 _09390_ (.A1(\core.decoded_imm_j[1] ),
    .A2(_03658_),
    .B1(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__nand3_2 _09391_ (.A(\core.decoded_imm_j[1] ),
    .B(_03658_),
    .C(_03674_),
    .Y(_03676_));
 sky130_fd_sc_hd__buf_1 _09392_ (.A(_02108_),
    .X(_03677_));
 sky130_fd_sc_hd__a32o_2 _09393_ (.A1(_03673_),
    .A2(_03675_),
    .A3(_03676_),
    .B1(_03670_),
    .B2(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__o221a_2 _09394_ (.A1(_03655_),
    .A2(\core.reg_next_pc[2] ),
    .B1(_03671_),
    .B2(_03678_),
    .C1(_03665_),
    .X(_00118_));
 sky130_fd_sc_hd__buf_1 _09395_ (.A(_02080_),
    .X(_03679_));
 sky130_fd_sc_hd__buf_1 _09396_ (.A(_03486_),
    .X(_03680_));
 sky130_fd_sc_hd__buf_1 _09397_ (.A(_02110_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_2 _09398_ (.A0(\core.reg_out[3] ),
    .A1(\core.alu_out_q[3] ),
    .S(\core.latched_stalu ),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_2 _09399_ (.A0(_03682_),
    .A1(\core.reg_next_pc[3] ),
    .S(_03199_),
    .X(_03683_));
 sky130_fd_sc_hd__or2_2 _09400_ (.A(_03681_),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__nand2_2 _09401_ (.A(\core.cpu_state[1] ),
    .B(\core.decoder_trigger ),
    .Y(_03685_));
 sky130_fd_sc_hd__buf_1 _09402_ (.A(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__nand2_2 _09403_ (.A(\core.decoded_imm_j[3] ),
    .B(_03683_),
    .Y(_03687_));
 sky130_fd_sc_hd__or2_2 _09404_ (.A(\core.decoded_imm_j[3] ),
    .B(_03683_),
    .X(_03688_));
 sky130_fd_sc_hd__nand2_2 _09405_ (.A(_03687_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__and2_2 _09406_ (.A(\core.decoded_imm_j[2] ),
    .B(_03670_),
    .X(_03690_));
 sky130_fd_sc_hd__a31oi_2 _09407_ (.A1(\core.decoded_imm_j[1] ),
    .A2(_03658_),
    .A3(_03674_),
    .B1(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_2 _09408_ (.A(_03689_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__buf_1 _09409_ (.A(\core.instr_jal ),
    .X(_03693_));
 sky130_fd_sc_hd__nor2_2 _09410_ (.A(_03670_),
    .B(_03683_),
    .Y(_03694_));
 sky130_fd_sc_hd__and2_2 _09411_ (.A(_03670_),
    .B(_03683_),
    .X(_03695_));
 sky130_fd_sc_hd__or3_2 _09412_ (.A(_03693_),
    .B(_03694_),
    .C(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__o21ai_2 _09413_ (.A1(_03666_),
    .A2(_03692_),
    .B1(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__buf_1 _09414_ (.A(\core.decoder_trigger ),
    .X(_03698_));
 sky130_fd_sc_hd__a22o_2 _09415_ (.A1(_03684_),
    .A2(_03686_),
    .B1(_03697_),
    .B2(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__o211a_2 _09416_ (.A1(_03679_),
    .A2(\core.reg_next_pc[3] ),
    .B1(_03680_),
    .C1(_03699_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_2 _09417_ (.A0(\core.reg_out[4] ),
    .A1(\core.alu_out_q[4] ),
    .S(\core.latched_stalu ),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_2 _09418_ (.A0(_03700_),
    .A1(\core.reg_next_pc[4] ),
    .S(_03199_),
    .X(_03701_));
 sky130_fd_sc_hd__nor2_2 _09419_ (.A(_03695_),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__a31o_2 _09420_ (.A1(_03670_),
    .A2(_03683_),
    .A3(_03701_),
    .B1(\core.instr_jal ),
    .X(_03703_));
 sky130_fd_sc_hd__and2_2 _09421_ (.A(\core.decoded_imm_j[4] ),
    .B(_03701_),
    .X(_03704_));
 sky130_fd_sc_hd__nor2_2 _09422_ (.A(\core.decoded_imm_j[4] ),
    .B(_03701_),
    .Y(_03705_));
 sky130_fd_sc_hd__nor2_2 _09423_ (.A(_03704_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__nor2_2 _09424_ (.A(\core.decoded_imm_j[3] ),
    .B(_03683_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ai_2 _09425_ (.A1(_03707_),
    .A2(_03691_),
    .B1(_03687_),
    .Y(_03708_));
 sky130_fd_sc_hd__xor2_2 _09426_ (.A(_03706_),
    .B(_03708_),
    .X(_03709_));
 sky130_fd_sc_hd__a2bb2o_2 _09427_ (.A1_N(_03702_),
    .A2_N(_03703_),
    .B1(_03709_),
    .B2(_02018_),
    .X(_03710_));
 sky130_fd_sc_hd__or2_2 _09428_ (.A(_03663_),
    .B(_03701_),
    .X(_03711_));
 sky130_fd_sc_hd__a22o_2 _09429_ (.A1(_03698_),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03686_),
    .X(_03712_));
 sky130_fd_sc_hd__o211a_2 _09430_ (.A1(_03679_),
    .A2(\core.reg_next_pc[4] ),
    .B1(_03680_),
    .C1(_03712_),
    .X(_00120_));
 sky130_fd_sc_hd__buf_1 _09431_ (.A(_02111_),
    .X(_03713_));
 sky130_fd_sc_hd__buf_1 _09432_ (.A(_03693_),
    .X(_03714_));
 sky130_fd_sc_hd__a21o_2 _09433_ (.A1(_03706_),
    .A2(_03708_),
    .B1(_03704_),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_2 _09434_ (.A0(\core.reg_out[5] ),
    .A1(\core.alu_out_q[5] ),
    .S(\core.latched_stalu ),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_2 _09435_ (.A0(_03716_),
    .A1(\core.reg_next_pc[5] ),
    .S(_03199_),
    .X(_03717_));
 sky130_fd_sc_hd__nor2_2 _09436_ (.A(\core.decoded_imm_j[5] ),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__and2_2 _09437_ (.A(\core.decoded_imm_j[5] ),
    .B(_03717_),
    .X(_03719_));
 sky130_fd_sc_hd__nor2_2 _09438_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__and2_2 _09439_ (.A(_03715_),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__inv_2 _09440_ (.A(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__or2_2 _09441_ (.A(_03715_),
    .B(_03720_),
    .X(_03723_));
 sky130_fd_sc_hd__and4_2 _09442_ (.A(_03670_),
    .B(_03683_),
    .C(_03701_),
    .D(_03717_),
    .X(_03724_));
 sky130_fd_sc_hd__o21ai_2 _09443_ (.A1(_03714_),
    .A2(_03724_),
    .B1(_03659_),
    .Y(_03725_));
 sky130_fd_sc_hd__a31o_2 _09444_ (.A1(_03714_),
    .A2(_03722_),
    .A3(_03723_),
    .B1(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__a21o_2 _09445_ (.A1(_03698_),
    .A2(_03703_),
    .B1(_03717_),
    .X(_03727_));
 sky130_fd_sc_hd__nor2_2 _09446_ (.A(\core.cpu_state[1] ),
    .B(_02048_),
    .Y(_03728_));
 sky130_fd_sc_hd__buf_1 _09447_ (.A(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a32o_2 _09448_ (.A1(_03713_),
    .A2(_03726_),
    .A3(_03727_),
    .B1(_03729_),
    .B2(\core.reg_next_pc[5] ),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_2 _09449_ (.A0(\core.reg_out[6] ),
    .A1(\core.alu_out_q[6] ),
    .S(_03656_),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_2 _09450_ (.A0(_03730_),
    .A1(\core.reg_next_pc[6] ),
    .S(_03200_),
    .X(_03731_));
 sky130_fd_sc_hd__nand2_2 _09451_ (.A(_03724_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__and2_2 _09452_ (.A(\core.decoded_imm_j[6] ),
    .B(_03731_),
    .X(_03733_));
 sky130_fd_sc_hd__or2_2 _09453_ (.A(\core.decoded_imm_j[6] ),
    .B(_03731_),
    .X(_03734_));
 sky130_fd_sc_hd__and2b_2 _09454_ (.A_N(_03733_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__o21ai_2 _09455_ (.A1(_03719_),
    .A2(_03721_),
    .B1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__o31a_2 _09456_ (.A1(_03719_),
    .A2(_03721_),
    .A3(_03735_),
    .B1(_03693_),
    .X(_03737_));
 sky130_fd_sc_hd__a221o_2 _09457_ (.A1(_03666_),
    .A2(_03732_),
    .B1(_03736_),
    .B2(_03737_),
    .C1(_03677_),
    .X(_03738_));
 sky130_fd_sc_hd__or2b_2 _09458_ (.A(_03731_),
    .B_N(_03725_),
    .X(_03739_));
 sky130_fd_sc_hd__a32o_2 _09459_ (.A1(_03713_),
    .A2(_03738_),
    .A3(_03739_),
    .B1(_03729_),
    .B2(\core.reg_next_pc[6] ),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_2 _09460_ (.A0(\core.reg_out[7] ),
    .A1(\core.alu_out_q[7] ),
    .S(_03656_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_2 _09461_ (.A0(_03740_),
    .A1(\core.reg_next_pc[7] ),
    .S(_03199_),
    .X(_03741_));
 sky130_fd_sc_hd__nor2_2 _09462_ (.A(\core.decoded_imm_j[7] ),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__and2_2 _09463_ (.A(\core.decoded_imm_j[7] ),
    .B(_03741_),
    .X(_03743_));
 sky130_fd_sc_hd__nor2_2 _09464_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__o31a_2 _09465_ (.A1(_03719_),
    .A2(_03721_),
    .A3(_03733_),
    .B1(_03734_),
    .X(_03745_));
 sky130_fd_sc_hd__xnor2_2 _09466_ (.A(_03744_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__nor2_2 _09467_ (.A(_03672_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__or2_2 _09468_ (.A(_03681_),
    .B(_03741_),
    .X(_03748_));
 sky130_fd_sc_hd__xnor2_2 _09469_ (.A(_03732_),
    .B(_03741_),
    .Y(_03749_));
 sky130_fd_sc_hd__a22o_2 _09470_ (.A1(_03685_),
    .A2(_03748_),
    .B1(_03749_),
    .B2(_02109_),
    .X(_03750_));
 sky130_fd_sc_hd__o221a_2 _09471_ (.A1(_03655_),
    .A2(\core.reg_next_pc[7] ),
    .B1(_03747_),
    .B2(_03750_),
    .C1(_03665_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_2 _09472_ (.A0(\core.reg_out[8] ),
    .A1(\core.alu_out_q[8] ),
    .S(_03656_),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_2 _09473_ (.A0(_03751_),
    .A1(\core.reg_next_pc[8] ),
    .S(_03199_),
    .X(_03752_));
 sky130_fd_sc_hd__a31oi_2 _09474_ (.A1(_03724_),
    .A2(_03731_),
    .A3(_03741_),
    .B1(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand4_2 _09475_ (.A(_03724_),
    .B(_03731_),
    .C(_03741_),
    .D(_03752_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_2 _09476_ (.A(_03666_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__or2_2 _09477_ (.A(\core.decoded_imm_j[8] ),
    .B(_03752_),
    .X(_03756_));
 sky130_fd_sc_hd__nand2_2 _09478_ (.A(\core.decoded_imm_j[8] ),
    .B(_03752_),
    .Y(_03757_));
 sky130_fd_sc_hd__and2_2 _09479_ (.A(_03756_),
    .B(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__a21o_2 _09480_ (.A1(_03744_),
    .A2(_03745_),
    .B1(_03743_),
    .X(_03759_));
 sky130_fd_sc_hd__xor2_2 _09481_ (.A(_03758_),
    .B(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__a2bb2o_2 _09482_ (.A1_N(_03753_),
    .A2_N(_03755_),
    .B1(_03760_),
    .B2(_02018_),
    .X(_03761_));
 sky130_fd_sc_hd__or2_2 _09483_ (.A(_03663_),
    .B(_03752_),
    .X(_03762_));
 sky130_fd_sc_hd__a22o_2 _09484_ (.A1(_03698_),
    .A2(_03761_),
    .B1(_03762_),
    .B2(_03686_),
    .X(_03763_));
 sky130_fd_sc_hd__o211a_2 _09485_ (.A1(_03679_),
    .A2(\core.reg_next_pc[8] ),
    .B1(_03680_),
    .C1(_03763_),
    .X(_00124_));
 sky130_fd_sc_hd__and4_2 _09486_ (.A(_03715_),
    .B(_03720_),
    .C(_03744_),
    .D(_03758_),
    .X(_03764_));
 sky130_fd_sc_hd__a31o_2 _09487_ (.A1(\core.decoded_imm_j[5] ),
    .A2(_03717_),
    .A3(_03734_),
    .B1(_03733_),
    .X(_03765_));
 sky130_fd_sc_hd__and3_2 _09488_ (.A(_03744_),
    .B(_03758_),
    .C(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__inv_2 _09489_ (.A(_03757_),
    .Y(_03767_));
 sky130_fd_sc_hd__a31o_2 _09490_ (.A1(\core.decoded_imm_j[7] ),
    .A2(_03741_),
    .A3(_03756_),
    .B1(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a211o_2 _09491_ (.A1(_03735_),
    .A2(_03764_),
    .B1(_03766_),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_2 _09492_ (.A0(\core.reg_out[9] ),
    .A1(\core.alu_out_q[9] ),
    .S(\core.latched_stalu ),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_2 _09493_ (.A0(_03770_),
    .A1(\core.reg_next_pc[9] ),
    .S(_03199_),
    .X(_03771_));
 sky130_fd_sc_hd__xor2_2 _09494_ (.A(\core.decoded_imm_j[9] ),
    .B(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__nand2_2 _09495_ (.A(_03769_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__or2_2 _09496_ (.A(_03769_),
    .B(_03772_),
    .X(_03774_));
 sky130_fd_sc_hd__inv_2 _09497_ (.A(_03771_),
    .Y(_03775_));
 sky130_fd_sc_hd__o21ai_2 _09498_ (.A1(_03754_),
    .A2(_03775_),
    .B1(_03666_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand2_2 _09499_ (.A(\core.decoder_trigger ),
    .B(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__a31o_2 _09500_ (.A1(_03714_),
    .A2(_03773_),
    .A3(_03774_),
    .B1(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__a21o_2 _09501_ (.A1(_03659_),
    .A2(_03755_),
    .B1(_03771_),
    .X(_03779_));
 sky130_fd_sc_hd__a32o_2 _09502_ (.A1(_03713_),
    .A2(_03778_),
    .A3(_03779_),
    .B1(_03729_),
    .B2(\core.reg_next_pc[9] ),
    .X(_00125_));
 sky130_fd_sc_hd__buf_1 _09503_ (.A(_03728_),
    .X(_03780_));
 sky130_fd_sc_hd__mux2_2 _09504_ (.A0(\core.reg_out[10] ),
    .A1(\core.alu_out_q[10] ),
    .S(_03656_),
    .X(_03781_));
 sky130_fd_sc_hd__mux2_2 _09505_ (.A0(_03781_),
    .A1(\core.reg_next_pc[10] ),
    .S(_03200_),
    .X(_03782_));
 sky130_fd_sc_hd__or2_2 _09506_ (.A(\core.decoded_imm_j[10] ),
    .B(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__inv_2 _09507_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__and2_2 _09508_ (.A(\core.decoded_imm_j[10] ),
    .B(_03782_),
    .X(_03785_));
 sky130_fd_sc_hd__nor2_2 _09509_ (.A(_03784_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__a21bo_2 _09510_ (.A1(\core.decoded_imm_j[9] ),
    .A2(_03771_),
    .B1_N(_03773_),
    .X(_03787_));
 sky130_fd_sc_hd__xnor2_2 _09511_ (.A(_03786_),
    .B(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__inv_2 _09512_ (.A(_03782_),
    .Y(_03789_));
 sky130_fd_sc_hd__and3b_2 _09513_ (.A_N(_03754_),
    .B(_03771_),
    .C(_03782_),
    .X(_03790_));
 sky130_fd_sc_hd__nand2_2 _09514_ (.A(_02079_),
    .B(_02024_),
    .Y(_03791_));
 sky130_fd_sc_hd__a221o_2 _09515_ (.A1(_03777_),
    .A2(_03789_),
    .B1(_03790_),
    .B2(_02109_),
    .C1(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__a21oi_2 _09516_ (.A1(_03673_),
    .A2(_03788_),
    .B1(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__a21o_2 _09517_ (.A1(\core.reg_next_pc[10] ),
    .A2(_03780_),
    .B1(_03793_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_2 _09518_ (.A0(\core.reg_out[11] ),
    .A1(\core.alu_out_q[11] ),
    .S(_03656_),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_2 _09519_ (.A0(_03794_),
    .A1(\core.reg_next_pc[11] ),
    .S(_03200_),
    .X(_03795_));
 sky130_fd_sc_hd__nor2_2 _09520_ (.A(\core.decoded_imm_j[11] ),
    .B(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__and2_2 _09521_ (.A(\core.decoded_imm_j[11] ),
    .B(_03795_),
    .X(_03797_));
 sky130_fd_sc_hd__nor2_2 _09522_ (.A(_03796_),
    .B(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__o21a_2 _09523_ (.A1(_03785_),
    .A2(_03787_),
    .B1(_03783_),
    .X(_03799_));
 sky130_fd_sc_hd__o21ai_2 _09524_ (.A1(_03798_),
    .A2(_03799_),
    .B1(_03673_),
    .Y(_03800_));
 sky130_fd_sc_hd__a21oi_2 _09525_ (.A1(_03798_),
    .A2(_03799_),
    .B1(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__or2_2 _09526_ (.A(_03790_),
    .B(_03795_),
    .X(_03802_));
 sky130_fd_sc_hd__or4bb_2 _09527_ (.A(_03754_),
    .B(_03775_),
    .C_N(_03782_),
    .D_N(_03795_),
    .X(_03803_));
 sky130_fd_sc_hd__or2_2 _09528_ (.A(_03681_),
    .B(_03795_),
    .X(_03804_));
 sky130_fd_sc_hd__a32o_2 _09529_ (.A1(_02109_),
    .A2(_03802_),
    .A3(_03803_),
    .B1(_03686_),
    .B2(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__o221a_2 _09530_ (.A1(_03655_),
    .A2(\core.reg_next_pc[11] ),
    .B1(_03801_),
    .B2(_03805_),
    .C1(_03665_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_2 _09531_ (.A0(\core.reg_out[12] ),
    .A1(\core.alu_out_q[12] ),
    .S(_03656_),
    .X(_03806_));
 sky130_fd_sc_hd__and3_2 _09532_ (.A(\core.latched_store ),
    .B(\core.latched_branch ),
    .C(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a21oi_2 _09533_ (.A1(\core.reg_next_pc[12] ),
    .A2(_03201_),
    .B1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_2 _09534_ (.A(_03803_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__nor2_2 _09535_ (.A(_03803_),
    .B(_03808_),
    .Y(_03810_));
 sky130_fd_sc_hd__nor2_2 _09536_ (.A(_03693_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__mux2_2 _09537_ (.A0(_03806_),
    .A1(\core.reg_next_pc[12] ),
    .S(_03200_),
    .X(_03812_));
 sky130_fd_sc_hd__xor2_2 _09538_ (.A(\core.decoded_imm_j[12] ),
    .B(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__a21oi_2 _09539_ (.A1(_03798_),
    .A2(_03799_),
    .B1(_03797_),
    .Y(_03814_));
 sky130_fd_sc_hd__xnor2_2 _09540_ (.A(_03813_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__a22o_2 _09541_ (.A1(_03809_),
    .A2(_03811_),
    .B1(_03815_),
    .B2(_02018_),
    .X(_03816_));
 sky130_fd_sc_hd__or2_2 _09542_ (.A(_03663_),
    .B(_03812_),
    .X(_03817_));
 sky130_fd_sc_hd__a22o_2 _09543_ (.A1(_03698_),
    .A2(_03816_),
    .B1(_03817_),
    .B2(_03686_),
    .X(_03818_));
 sky130_fd_sc_hd__o211a_2 _09544_ (.A1(_03679_),
    .A2(\core.reg_next_pc[12] ),
    .B1(_03680_),
    .C1(_03818_),
    .X(_00128_));
 sky130_fd_sc_hd__a31o_2 _09545_ (.A1(\core.decoded_imm_j[9] ),
    .A2(_03771_),
    .A3(_03783_),
    .B1(_03785_),
    .X(_03819_));
 sky130_fd_sc_hd__o211a_2 _09546_ (.A1(\core.decoded_imm_j[12] ),
    .A2(_03812_),
    .B1(_03795_),
    .C1(\core.decoded_imm_j[11] ),
    .X(_03820_));
 sky130_fd_sc_hd__a21o_2 _09547_ (.A1(\core.decoded_imm_j[12] ),
    .A2(_03812_),
    .B1(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__a31o_2 _09548_ (.A1(_03798_),
    .A2(_03813_),
    .A3(_03819_),
    .B1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__and4_2 _09549_ (.A(_03772_),
    .B(_03786_),
    .C(_03798_),
    .D(_03813_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_2 _09550_ (.A(_03769_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__mux2_2 _09551_ (.A0(\core.reg_out[13] ),
    .A1(\core.alu_out_q[13] ),
    .S(_03656_),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_2 _09552_ (.A0(_03825_),
    .A1(\core.reg_next_pc[13] ),
    .S(_03200_),
    .X(_03826_));
 sky130_fd_sc_hd__buf_1 _09553_ (.A(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__xor2_2 _09554_ (.A(\core.decoded_imm_j[13] ),
    .B(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__o21a_2 _09555_ (.A1(_03822_),
    .A2(_03824_),
    .B1(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__o31ai_2 _09556_ (.A1(_03828_),
    .A2(_03822_),
    .A3(_03824_),
    .B1(_03714_),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_2 _09557_ (.A(_03810_),
    .B(_03827_),
    .Y(_03831_));
 sky130_fd_sc_hd__a21oi_2 _09558_ (.A1(_03666_),
    .A2(_03831_),
    .B1(_02108_),
    .Y(_03832_));
 sky130_fd_sc_hd__o21ai_2 _09559_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__o21a_2 _09560_ (.A1(_03693_),
    .A2(_03810_),
    .B1(\core.decoder_trigger ),
    .X(_03834_));
 sky130_fd_sc_hd__or2_2 _09561_ (.A(_03827_),
    .B(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__a32o_2 _09562_ (.A1(_03713_),
    .A2(_03833_),
    .A3(_03835_),
    .B1(_03729_),
    .B2(\core.reg_next_pc[13] ),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_2 _09563_ (.A0(\core.reg_out[14] ),
    .A1(\core.alu_out_q[14] ),
    .S(_03656_),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_2 _09564_ (.A0(_03836_),
    .A1(\core.reg_next_pc[14] ),
    .S(_03200_),
    .X(_03837_));
 sky130_fd_sc_hd__nand2_2 _09565_ (.A(\core.decoded_imm_j[14] ),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__or2_2 _09566_ (.A(\core.decoded_imm_j[14] ),
    .B(_03837_),
    .X(_03839_));
 sky130_fd_sc_hd__a21oi_2 _09567_ (.A1(\core.decoded_imm_j[13] ),
    .A2(_03827_),
    .B1(_03829_),
    .Y(_03840_));
 sky130_fd_sc_hd__a21oi_2 _09568_ (.A1(_03838_),
    .A2(_03839_),
    .B1(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__a31o_2 _09569_ (.A1(_03838_),
    .A2(_03839_),
    .A3(_03840_),
    .B1(_03672_),
    .X(_03842_));
 sky130_fd_sc_hd__nor2_2 _09570_ (.A(_03841_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__or4bb_2 _09571_ (.A(_03803_),
    .B(_03808_),
    .C_N(_03827_),
    .D_N(_03837_),
    .X(_03844_));
 sky130_fd_sc_hd__o221ai_2 _09572_ (.A1(_03832_),
    .A2(_03837_),
    .B1(_03844_),
    .B2(_03667_),
    .C1(_02111_),
    .Y(_03845_));
 sky130_fd_sc_hd__a2bb2o_2 _09573_ (.A1_N(_03843_),
    .A2_N(_03845_),
    .B1(\core.reg_next_pc[14] ),
    .B2(_03780_),
    .X(_00130_));
 sky130_fd_sc_hd__buf_1 _09574_ (.A(_03656_),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_2 _09575_ (.A0(\core.reg_out[15] ),
    .A1(\core.alu_out_q[15] ),
    .S(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__mux2_2 _09576_ (.A0(_03847_),
    .A1(\core.reg_next_pc[15] ),
    .S(_03201_),
    .X(_03848_));
 sky130_fd_sc_hd__or2_2 _09577_ (.A(\core.decoded_imm_j[15] ),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_2 _09578_ (.A(\core.decoded_imm_j[15] ),
    .B(_03848_),
    .Y(_03850_));
 sky130_fd_sc_hd__and2_2 _09579_ (.A(_03849_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__inv_2 _09580_ (.A(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__a21bo_2 _09581_ (.A1(_03838_),
    .A2(_03840_),
    .B1_N(_03839_),
    .X(_03853_));
 sky130_fd_sc_hd__a21o_2 _09582_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03672_),
    .X(_03854_));
 sky130_fd_sc_hd__o21ba_2 _09583_ (.A1(_03852_),
    .A2(_03853_),
    .B1_N(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__or2_2 _09584_ (.A(_03681_),
    .B(_03848_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _09585_ (.A(_03848_),
    .Y(_03857_));
 sky130_fd_sc_hd__nand2_2 _09586_ (.A(_03844_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__nor2_2 _09587_ (.A(_03844_),
    .B(_03857_),
    .Y(_03859_));
 sky130_fd_sc_hd__nor2_2 _09588_ (.A(_03667_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__a22o_2 _09589_ (.A1(_03685_),
    .A2(_03856_),
    .B1(_03858_),
    .B2(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__o221a_2 _09590_ (.A1(_03655_),
    .A2(\core.reg_next_pc[15] ),
    .B1(_03855_),
    .B2(_03861_),
    .C1(_03665_),
    .X(_00131_));
 sky130_fd_sc_hd__buf_1 _09591_ (.A(_03846_),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_2 _09592_ (.A0(\core.reg_out[16] ),
    .A1(\core.alu_out_q[16] ),
    .S(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_2 _09593_ (.A0(_03863_),
    .A1(\core.reg_next_pc[16] ),
    .S(_03201_),
    .X(_03864_));
 sky130_fd_sc_hd__nor2_2 _09594_ (.A(_03859_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21o_2 _09595_ (.A1(_03859_),
    .A2(_03864_),
    .B1(_03693_),
    .X(_03866_));
 sky130_fd_sc_hd__xor2_2 _09596_ (.A(\core.decoded_imm_j[16] ),
    .B(_03864_),
    .X(_03867_));
 sky130_fd_sc_hd__o21ai_2 _09597_ (.A1(_03852_),
    .A2(_03853_),
    .B1(_03850_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_2 _09598_ (.A(_03867_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o22a_2 _09599_ (.A1(_03865_),
    .A2(_03866_),
    .B1(_03869_),
    .B2(_03666_),
    .X(_03870_));
 sky130_fd_sc_hd__nor2_2 _09600_ (.A(_03677_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__a21o_2 _09601_ (.A1(_03677_),
    .A2(_03864_),
    .B1(_03663_),
    .X(_03872_));
 sky130_fd_sc_hd__o221a_2 _09602_ (.A1(_03655_),
    .A2(\core.reg_next_pc[16] ),
    .B1(_03871_),
    .B2(_03872_),
    .C1(_03665_),
    .X(_00132_));
 sky130_fd_sc_hd__and3_2 _09603_ (.A(_03828_),
    .B(_03838_),
    .C(_03839_),
    .X(_03873_));
 sky130_fd_sc_hd__and3_2 _09604_ (.A(_03851_),
    .B(_03867_),
    .C(_03873_),
    .X(_03874_));
 sky130_fd_sc_hd__o21a_2 _09605_ (.A1(\core.decoded_imm_j[13] ),
    .A2(_03827_),
    .B1(_03822_),
    .X(_03875_));
 sky130_fd_sc_hd__a22o_2 _09606_ (.A1(\core.decoded_imm_j[13] ),
    .A2(_03827_),
    .B1(_03837_),
    .B2(\core.decoded_imm_j[14] ),
    .X(_03876_));
 sky130_fd_sc_hd__o211a_2 _09607_ (.A1(_03875_),
    .A2(_03876_),
    .B1(_03839_),
    .C1(_03849_),
    .X(_03877_));
 sky130_fd_sc_hd__a22o_2 _09608_ (.A1(\core.decoded_imm_j[15] ),
    .A2(_03848_),
    .B1(_03864_),
    .B2(\core.decoded_imm_j[16] ),
    .X(_03878_));
 sky130_fd_sc_hd__o22a_2 _09609_ (.A1(\core.decoded_imm_j[16] ),
    .A2(_03864_),
    .B1(_03877_),
    .B2(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__a31o_2 _09610_ (.A1(_03769_),
    .A2(_03823_),
    .A3(_03874_),
    .B1(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_2 _09611_ (.A0(\core.reg_out[17] ),
    .A1(\core.alu_out_q[17] ),
    .S(_03846_),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_2 _09612_ (.A0(_03881_),
    .A1(\core.reg_next_pc[17] ),
    .S(_03201_),
    .X(_03882_));
 sky130_fd_sc_hd__nor2_2 _09613_ (.A(\core.decoded_imm_j[17] ),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__and2_2 _09614_ (.A(\core.decoded_imm_j[17] ),
    .B(_03882_),
    .X(_03884_));
 sky130_fd_sc_hd__nor2_2 _09615_ (.A(_03883_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_2 _09616_ (.A(_03880_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__or2_2 _09617_ (.A(_03880_),
    .B(_03885_),
    .X(_03887_));
 sky130_fd_sc_hd__and4b_2 _09618_ (.A_N(_03844_),
    .B(_03848_),
    .C(_03864_),
    .D(_03882_),
    .X(_03888_));
 sky130_fd_sc_hd__o21ai_2 _09619_ (.A1(_03714_),
    .A2(_03888_),
    .B1(_03659_),
    .Y(_03889_));
 sky130_fd_sc_hd__a31o_2 _09620_ (.A1(_03714_),
    .A2(_03886_),
    .A3(_03887_),
    .B1(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__a21o_2 _09621_ (.A1(_03659_),
    .A2(_03866_),
    .B1(_03882_),
    .X(_03891_));
 sky130_fd_sc_hd__a32o_2 _09622_ (.A1(_03713_),
    .A2(_03890_),
    .A3(_03891_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[17] ),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_2 _09623_ (.A0(\core.reg_out[18] ),
    .A1(\core.alu_out_q[18] ),
    .S(_03846_),
    .X(_03892_));
 sky130_fd_sc_hd__mux2_2 _09624_ (.A0(_03892_),
    .A1(\core.reg_next_pc[18] ),
    .S(_03201_),
    .X(_03893_));
 sky130_fd_sc_hd__or2b_2 _09625_ (.A(_03893_),
    .B_N(_03889_),
    .X(_03894_));
 sky130_fd_sc_hd__and2_2 _09626_ (.A(\core.decoded_imm_j[18] ),
    .B(_03893_),
    .X(_03895_));
 sky130_fd_sc_hd__or2_2 _09627_ (.A(\core.decoded_imm_j[18] ),
    .B(_03893_),
    .X(_03896_));
 sky130_fd_sc_hd__and2b_2 _09628_ (.A_N(_03895_),
    .B(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a21o_2 _09629_ (.A1(_03880_),
    .A2(_03885_),
    .B1(_03884_),
    .X(_03898_));
 sky130_fd_sc_hd__xor2_2 _09630_ (.A(_03897_),
    .B(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_2 _09631_ (.A(_03888_),
    .B(_03893_),
    .Y(_03900_));
 sky130_fd_sc_hd__o22a_2 _09632_ (.A1(_03672_),
    .A2(_03899_),
    .B1(_03900_),
    .B2(_03667_),
    .X(_03901_));
 sky130_fd_sc_hd__a32o_2 _09633_ (.A1(_03713_),
    .A2(_03894_),
    .A3(_03901_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[18] ),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_2 _09634_ (.A0(\core.reg_out[19] ),
    .A1(\core.alu_out_q[19] ),
    .S(_03846_),
    .X(_03902_));
 sky130_fd_sc_hd__and3_2 _09635_ (.A(\core.latched_store ),
    .B(\core.latched_branch ),
    .C(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a21oi_2 _09636_ (.A1(\core.reg_next_pc[19] ),
    .A2(_03201_),
    .B1(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__xnor2_2 _09637_ (.A(\core.decoded_imm_j[19] ),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__o21a_2 _09638_ (.A1(_03895_),
    .A2(_03898_),
    .B1(_03896_),
    .X(_03906_));
 sky130_fd_sc_hd__and2_2 _09639_ (.A(_03905_),
    .B(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__nor2_2 _09640_ (.A(_03672_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__o21a_2 _09641_ (.A1(_03905_),
    .A2(_03906_),
    .B1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_2 _09642_ (.A(_02079_),
    .B(_03904_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_2 _09643_ (.A(_03900_),
    .B(_03904_),
    .Y(_03911_));
 sky130_fd_sc_hd__nor2_2 _09644_ (.A(_03900_),
    .B(_03904_),
    .Y(_03912_));
 sky130_fd_sc_hd__nor2_2 _09645_ (.A(_03667_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__a22o_2 _09646_ (.A1(_03685_),
    .A2(_03910_),
    .B1(_03911_),
    .B2(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__o221a_2 _09647_ (.A1(_03655_),
    .A2(\core.reg_next_pc[19] ),
    .B1(_03909_),
    .B2(_03914_),
    .C1(_03680_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_1 _09648_ (.A(_02082_),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_2 _09649_ (.A0(\core.reg_out[20] ),
    .A1(\core.alu_out_q[20] ),
    .S(_03846_),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_2 _09650_ (.A0(_03916_),
    .A1(\core.reg_next_pc[20] ),
    .S(_03201_),
    .X(_03917_));
 sky130_fd_sc_hd__nor2_2 _09651_ (.A(_03912_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21o_2 _09652_ (.A1(_03912_),
    .A2(_03917_),
    .B1(\core.instr_jal ),
    .X(_03919_));
 sky130_fd_sc_hd__buf_1 _09653_ (.A(\core.decoded_imm_j[20] ),
    .X(_03920_));
 sky130_fd_sc_hd__xor2_2 _09654_ (.A(_03920_),
    .B(_03917_),
    .X(_03921_));
 sky130_fd_sc_hd__inv_2 _09655_ (.A(_03904_),
    .Y(_03922_));
 sky130_fd_sc_hd__a21oi_2 _09656_ (.A1(\core.decoded_imm_j[19] ),
    .A2(_03922_),
    .B1(_03907_),
    .Y(_03923_));
 sky130_fd_sc_hd__xnor2_2 _09657_ (.A(_03921_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__a2bb2o_2 _09658_ (.A1_N(_03918_),
    .A2_N(_03919_),
    .B1(_02018_),
    .B2(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__or2_2 _09659_ (.A(_03681_),
    .B(_03917_),
    .X(_03926_));
 sky130_fd_sc_hd__a22o_2 _09660_ (.A1(_03698_),
    .A2(_03925_),
    .B1(_03926_),
    .B2(_03686_),
    .X(_03927_));
 sky130_fd_sc_hd__o211a_2 _09661_ (.A1(_03679_),
    .A2(\core.reg_next_pc[20] ),
    .B1(_03915_),
    .C1(_03927_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_2 _09662_ (.A0(\core.reg_out[21] ),
    .A1(\core.alu_out_q[21] ),
    .S(_03846_),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_2 _09663_ (.A0(_03928_),
    .A1(\core.reg_next_pc[21] ),
    .S(_03200_),
    .X(_03929_));
 sky130_fd_sc_hd__a21o_2 _09664_ (.A1(_03659_),
    .A2(_03919_),
    .B1(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_2 _09665_ (.A(_03920_),
    .B(_03929_),
    .Y(_03931_));
 sky130_fd_sc_hd__or2_2 _09666_ (.A(_03920_),
    .B(_03929_),
    .X(_03932_));
 sky130_fd_sc_hd__and2_2 _09667_ (.A(_03931_),
    .B(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__and2_2 _09668_ (.A(_03905_),
    .B(_03921_),
    .X(_03934_));
 sky130_fd_sc_hd__and3_2 _09669_ (.A(_03885_),
    .B(_03897_),
    .C(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_1 _09670_ (.A(_03920_),
    .X(_03936_));
 sky130_fd_sc_hd__a21o_2 _09671_ (.A1(_03884_),
    .A2(_03896_),
    .B1(_03895_),
    .X(_03937_));
 sky130_fd_sc_hd__o211a_2 _09672_ (.A1(_03936_),
    .A2(_03917_),
    .B1(_03922_),
    .C1(\core.decoded_imm_j[19] ),
    .X(_03938_));
 sky130_fd_sc_hd__a221o_2 _09673_ (.A1(_03936_),
    .A2(_03917_),
    .B1(_03934_),
    .B2(_03937_),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a21oi_2 _09674_ (.A1(_03880_),
    .A2(_03935_),
    .B1(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__xnor2_2 _09675_ (.A(_03933_),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__or4bb_2 _09676_ (.A(_03900_),
    .B(_03904_),
    .C_N(_03917_),
    .D_N(_03929_),
    .X(_03942_));
 sky130_fd_sc_hd__o22a_2 _09677_ (.A1(_03672_),
    .A2(_03941_),
    .B1(_03942_),
    .B2(_03667_),
    .X(_03943_));
 sky130_fd_sc_hd__a32o_2 _09678_ (.A1(_02111_),
    .A2(_03930_),
    .A3(_03943_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[21] ),
    .X(_00137_));
 sky130_fd_sc_hd__or2b_2 _09679_ (.A(_03940_),
    .B_N(_03933_),
    .X(_03944_));
 sky130_fd_sc_hd__mux2_2 _09680_ (.A0(\core.reg_out[22] ),
    .A1(\core.alu_out_q[22] ),
    .S(_03846_),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_2 _09681_ (.A0(_03945_),
    .A1(\core.reg_next_pc[22] ),
    .S(_03201_),
    .X(_03946_));
 sky130_fd_sc_hd__xnor2_2 _09682_ (.A(_03920_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__a21oi_2 _09683_ (.A1(_03931_),
    .A2(_03944_),
    .B1(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a31o_2 _09684_ (.A1(_03931_),
    .A2(_03944_),
    .A3(_03947_),
    .B1(_03666_),
    .X(_03949_));
 sky130_fd_sc_hd__or2_2 _09685_ (.A(_03948_),
    .B(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__and2b_2 _09686_ (.A_N(_03946_),
    .B(_03942_),
    .X(_03951_));
 sky130_fd_sc_hd__and2b_2 _09687_ (.A_N(_03942_),
    .B(_03946_),
    .X(_03952_));
 sky130_fd_sc_hd__or3_2 _09688_ (.A(_02018_),
    .B(_03951_),
    .C(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__a21oi_2 _09689_ (.A1(_03950_),
    .A2(_03953_),
    .B1(_03677_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21o_2 _09690_ (.A1(_03677_),
    .A2(_03946_),
    .B1(_03663_),
    .X(_03955_));
 sky130_fd_sc_hd__o221a_2 _09691_ (.A1(_03655_),
    .A2(\core.reg_next_pc[22] ),
    .B1(_03954_),
    .B2(_03955_),
    .C1(_03680_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_2 _09692_ (.A0(\core.reg_out[23] ),
    .A1(\core.alu_out_q[23] ),
    .S(_03846_),
    .X(_03956_));
 sky130_fd_sc_hd__mux2_2 _09693_ (.A0(_03956_),
    .A1(\core.reg_next_pc[23] ),
    .S(_03200_),
    .X(_03957_));
 sky130_fd_sc_hd__or2_2 _09694_ (.A(_03681_),
    .B(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__and2_2 _09695_ (.A(_03685_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__o21a_2 _09696_ (.A1(_03929_),
    .A2(_03946_),
    .B1(_03936_),
    .X(_03960_));
 sky130_fd_sc_hd__nor2_2 _09697_ (.A(_03944_),
    .B(_03947_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand2_2 _09698_ (.A(_03920_),
    .B(_03957_),
    .Y(_03962_));
 sky130_fd_sc_hd__or2_2 _09699_ (.A(_03920_),
    .B(_03957_),
    .X(_03963_));
 sky130_fd_sc_hd__and2_2 _09700_ (.A(_03962_),
    .B(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__o21ai_2 _09701_ (.A1(_03960_),
    .A2(_03961_),
    .B1(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__or3_2 _09702_ (.A(_03964_),
    .B(_03960_),
    .C(_03961_),
    .X(_03966_));
 sky130_fd_sc_hd__and2_2 _09703_ (.A(_03952_),
    .B(_03957_),
    .X(_03967_));
 sky130_fd_sc_hd__nor2_2 _09704_ (.A(_03667_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__o21a_2 _09705_ (.A1(_03952_),
    .A2(_03957_),
    .B1(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__a31o_2 _09706_ (.A1(_03673_),
    .A2(_03965_),
    .A3(_03966_),
    .B1(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__o221a_2 _09707_ (.A1(_02080_),
    .A2(\core.reg_next_pc[23] ),
    .B1(_03959_),
    .B2(_03970_),
    .C1(_03680_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_2 _09708_ (.A0(\core.reg_out[24] ),
    .A1(\core.alu_out_q[24] ),
    .S(_03846_),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_2 _09709_ (.A0(_03971_),
    .A1(\core.reg_next_pc[24] ),
    .S(_03201_),
    .X(_03972_));
 sky130_fd_sc_hd__xnor2_2 _09710_ (.A(_03920_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__a21oi_2 _09711_ (.A1(_03962_),
    .A2(_03965_),
    .B1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__a31o_2 _09712_ (.A1(_03962_),
    .A2(_03965_),
    .A3(_03973_),
    .B1(_03666_),
    .X(_03975_));
 sky130_fd_sc_hd__nor2_2 _09713_ (.A(_03974_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__a21oi_2 _09714_ (.A1(_03967_),
    .A2(_03972_),
    .B1(_03693_),
    .Y(_03977_));
 sky130_fd_sc_hd__o21a_2 _09715_ (.A1(_03967_),
    .A2(_03972_),
    .B1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__o21a_2 _09716_ (.A1(_03976_),
    .A2(_03978_),
    .B1(_03698_),
    .X(_03979_));
 sky130_fd_sc_hd__a21o_2 _09717_ (.A1(_03677_),
    .A2(_03972_),
    .B1(_03663_),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_2 _09718_ (.A1(_02080_),
    .A2(\core.reg_next_pc[24] ),
    .B1(_03979_),
    .B2(_03980_),
    .C1(_03680_),
    .X(_00140_));
 sky130_fd_sc_hd__inv_2 _09719_ (.A(_03947_),
    .Y(_03981_));
 sky130_fd_sc_hd__inv_2 _09720_ (.A(_03973_),
    .Y(_03982_));
 sky130_fd_sc_hd__and4_2 _09721_ (.A(_03933_),
    .B(_03981_),
    .C(_03964_),
    .D(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__and4_2 _09722_ (.A(_03885_),
    .B(_03897_),
    .C(_03934_),
    .D(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__o21a_2 _09723_ (.A1(_03957_),
    .A2(_03972_),
    .B1(_03936_),
    .X(_03985_));
 sky130_fd_sc_hd__a211o_2 _09724_ (.A1(_03939_),
    .A2(_03983_),
    .B1(_03985_),
    .C1(_03960_),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_2 _09725_ (.A1(_03880_),
    .A2(_03984_),
    .B1(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__mux2_2 _09726_ (.A0(\core.reg_out[25] ),
    .A1(\core.alu_out_q[25] ),
    .S(_03862_),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_2 _09727_ (.A0(_03988_),
    .A1(\core.reg_next_pc[25] ),
    .S(_03202_),
    .X(_03989_));
 sky130_fd_sc_hd__xor2_2 _09728_ (.A(_03936_),
    .B(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__or2b_2 _09729_ (.A(_03987_),
    .B_N(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__or2b_2 _09730_ (.A(_03990_),
    .B_N(_03987_),
    .X(_03992_));
 sky130_fd_sc_hd__and3_2 _09731_ (.A(_03967_),
    .B(_03972_),
    .C(_03989_),
    .X(_03993_));
 sky130_fd_sc_hd__o21ai_2 _09732_ (.A1(_03714_),
    .A2(_03993_),
    .B1(_03659_),
    .Y(_03994_));
 sky130_fd_sc_hd__a31o_2 _09733_ (.A1(_03714_),
    .A2(_03991_),
    .A3(_03992_),
    .B1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__o21bai_2 _09734_ (.A1(_03677_),
    .A2(_03977_),
    .B1_N(_03989_),
    .Y(_03996_));
 sky130_fd_sc_hd__a32o_2 _09735_ (.A1(_02111_),
    .A2(_03995_),
    .A3(_03996_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[25] ),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_2 _09736_ (.A0(\core.reg_out[26] ),
    .A1(\core.alu_out_q[26] ),
    .S(_03862_),
    .X(_03997_));
 sky130_fd_sc_hd__mux2_2 _09737_ (.A0(_03997_),
    .A1(\core.reg_next_pc[26] ),
    .S(_03202_),
    .X(_03998_));
 sky130_fd_sc_hd__xor2_2 _09738_ (.A(_03936_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__buf_1 _09739_ (.A(_03936_),
    .X(_04000_));
 sky130_fd_sc_hd__a21bo_2 _09740_ (.A1(_04000_),
    .A2(_03989_),
    .B1_N(_03991_),
    .X(_04001_));
 sky130_fd_sc_hd__xor2_2 _09741_ (.A(_03999_),
    .B(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__a21oi_2 _09742_ (.A1(_03993_),
    .A2(_03998_),
    .B1(_03693_),
    .Y(_04003_));
 sky130_fd_sc_hd__or2_2 _09743_ (.A(_03993_),
    .B(_03998_),
    .X(_04004_));
 sky130_fd_sc_hd__a22o_2 _09744_ (.A1(_02018_),
    .A2(_04002_),
    .B1(_04003_),
    .B2(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__or2_2 _09745_ (.A(_03681_),
    .B(_03998_),
    .X(_04006_));
 sky130_fd_sc_hd__a22o_2 _09746_ (.A1(_03698_),
    .A2(_04005_),
    .B1(_04006_),
    .B2(_03686_),
    .X(_04007_));
 sky130_fd_sc_hd__o211a_2 _09747_ (.A1(_03679_),
    .A2(\core.reg_next_pc[26] ),
    .B1(_03915_),
    .C1(_04007_),
    .X(_00142_));
 sky130_fd_sc_hd__o21a_2 _09748_ (.A1(_03989_),
    .A2(_03998_),
    .B1(_03936_),
    .X(_04008_));
 sky130_fd_sc_hd__and2b_2 _09749_ (.A_N(_03991_),
    .B(_03999_),
    .X(_04009_));
 sky130_fd_sc_hd__mux2_2 _09750_ (.A0(\core.reg_out[27] ),
    .A1(\core.alu_out_q[27] ),
    .S(_03862_),
    .X(_04010_));
 sky130_fd_sc_hd__mux2_2 _09751_ (.A0(_04010_),
    .A1(\core.reg_next_pc[27] ),
    .S(_03202_),
    .X(_04011_));
 sky130_fd_sc_hd__xor2_2 _09752_ (.A(_03936_),
    .B(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__o21a_2 _09753_ (.A1(_04008_),
    .A2(_04009_),
    .B1(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__nor3_2 _09754_ (.A(_04012_),
    .B(_04008_),
    .C(_04009_),
    .Y(_04014_));
 sky130_fd_sc_hd__o21ai_2 _09755_ (.A1(_04013_),
    .A2(_04014_),
    .B1(_03673_),
    .Y(_04015_));
 sky130_fd_sc_hd__o21bai_2 _09756_ (.A1(_03677_),
    .A2(_04003_),
    .B1_N(_04011_),
    .Y(_04016_));
 sky130_fd_sc_hd__and3_2 _09757_ (.A(_03993_),
    .B(_03998_),
    .C(_04011_),
    .X(_04017_));
 sky130_fd_sc_hd__a21oi_2 _09758_ (.A1(_02109_),
    .A2(_04017_),
    .B1(_03791_),
    .Y(_04018_));
 sky130_fd_sc_hd__a32o_2 _09759_ (.A1(_04015_),
    .A2(_04016_),
    .A3(_04018_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[27] ),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_2 _09760_ (.A0(\core.reg_out[28] ),
    .A1(\core.alu_out_q[28] ),
    .S(_03862_),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_2 _09761_ (.A0(_04019_),
    .A1(\core.reg_next_pc[28] ),
    .S(_03202_),
    .X(_04020_));
 sky130_fd_sc_hd__nor2_2 _09762_ (.A(_04017_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21o_2 _09763_ (.A1(_04017_),
    .A2(_04020_),
    .B1(\core.instr_jal ),
    .X(_04022_));
 sky130_fd_sc_hd__xor2_2 _09764_ (.A(_03936_),
    .B(_04020_),
    .X(_04023_));
 sky130_fd_sc_hd__a21o_2 _09765_ (.A1(_04000_),
    .A2(_04011_),
    .B1(_04013_),
    .X(_04024_));
 sky130_fd_sc_hd__xor2_2 _09766_ (.A(_04023_),
    .B(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__a2bb2o_2 _09767_ (.A1_N(_04021_),
    .A2_N(_04022_),
    .B1(_02018_),
    .B2(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__or2_2 _09768_ (.A(_03681_),
    .B(_04020_),
    .X(_04027_));
 sky130_fd_sc_hd__a22o_2 _09769_ (.A1(_03698_),
    .A2(_04026_),
    .B1(_04027_),
    .B2(_03686_),
    .X(_04028_));
 sky130_fd_sc_hd__o211a_2 _09770_ (.A1(_03679_),
    .A2(\core.reg_next_pc[28] ),
    .B1(_03915_),
    .C1(_04028_),
    .X(_00144_));
 sky130_fd_sc_hd__o21a_2 _09771_ (.A1(_04011_),
    .A2(_04020_),
    .B1(_04000_),
    .X(_04029_));
 sky130_fd_sc_hd__a311o_2 _09772_ (.A1(_04012_),
    .A2(_04009_),
    .A3(_04023_),
    .B1(_04029_),
    .C1(_04008_),
    .X(_04030_));
 sky130_fd_sc_hd__mux2_2 _09773_ (.A0(\core.reg_out[29] ),
    .A1(\core.alu_out_q[29] ),
    .S(_03862_),
    .X(_04031_));
 sky130_fd_sc_hd__mux2_2 _09774_ (.A0(_04031_),
    .A1(\core.reg_next_pc[29] ),
    .S(_03202_),
    .X(_04032_));
 sky130_fd_sc_hd__and2_2 _09775_ (.A(_04000_),
    .B(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__or2_2 _09776_ (.A(_04000_),
    .B(_04032_),
    .X(_04034_));
 sky130_fd_sc_hd__or2b_2 _09777_ (.A(_04033_),
    .B_N(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__xnor2_2 _09778_ (.A(_04030_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__and3_2 _09779_ (.A(_04017_),
    .B(_04020_),
    .C(_04032_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_2 _09780_ (.A(_03714_),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__a211o_2 _09781_ (.A1(_03714_),
    .A2(_04036_),
    .B1(_04038_),
    .C1(_03677_),
    .X(_04039_));
 sky130_fd_sc_hd__a21o_2 _09782_ (.A1(_03659_),
    .A2(_04022_),
    .B1(_04032_),
    .X(_04040_));
 sky130_fd_sc_hd__a32o_2 _09783_ (.A1(_02111_),
    .A2(_04039_),
    .A3(_04040_),
    .B1(_03728_),
    .B2(\core.reg_next_pc[29] ),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_2 _09784_ (.A0(\core.reg_out[30] ),
    .A1(\core.alu_out_q[30] ),
    .S(_03862_),
    .X(_04041_));
 sky130_fd_sc_hd__mux2_2 _09785_ (.A0(_04041_),
    .A1(\core.reg_next_pc[30] ),
    .S(_03202_),
    .X(_04042_));
 sky130_fd_sc_hd__or2_2 _09786_ (.A(_04000_),
    .B(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__nand2_2 _09787_ (.A(_04000_),
    .B(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__a21o_2 _09788_ (.A1(_04030_),
    .A2(_04034_),
    .B1(_04033_),
    .X(_04045_));
 sky130_fd_sc_hd__a21oi_2 _09789_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__a31o_2 _09790_ (.A1(_04043_),
    .A2(_04044_),
    .A3(_04045_),
    .B1(_03672_),
    .X(_04047_));
 sky130_fd_sc_hd__nor2_2 _09791_ (.A(_04046_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__or2_2 _09792_ (.A(_04037_),
    .B(_04042_),
    .X(_04049_));
 sky130_fd_sc_hd__nand2_2 _09793_ (.A(_04037_),
    .B(_04042_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_2 _09794_ (.A(_03681_),
    .B(_04042_),
    .X(_04051_));
 sky130_fd_sc_hd__a32o_2 _09795_ (.A1(_02109_),
    .A2(_04049_),
    .A3(_04050_),
    .B1(_03686_),
    .B2(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__o221a_2 _09796_ (.A1(_02080_),
    .A2(\core.reg_next_pc[30] ),
    .B1(_04048_),
    .B2(_04052_),
    .C1(_03680_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_2 _09797_ (.A0(\core.reg_out[31] ),
    .A1(\core.alu_out_q[31] ),
    .S(_03862_),
    .X(_04053_));
 sky130_fd_sc_hd__mux2_2 _09798_ (.A0(_04053_),
    .A1(\core.reg_next_pc[31] ),
    .S(_03202_),
    .X(_04054_));
 sky130_fd_sc_hd__xnor2_2 _09799_ (.A(_04050_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__a21bo_2 _09800_ (.A1(_04043_),
    .A2(_04045_),
    .B1_N(_04044_),
    .X(_04056_));
 sky130_fd_sc_hd__xnor2_2 _09801_ (.A(_04000_),
    .B(_04054_),
    .Y(_04057_));
 sky130_fd_sc_hd__xnor2_2 _09802_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__mux2_2 _09803_ (.A0(_04055_),
    .A1(_04058_),
    .S(_03693_),
    .X(_04059_));
 sky130_fd_sc_hd__or2_2 _09804_ (.A(_03681_),
    .B(_04054_),
    .X(_04060_));
 sky130_fd_sc_hd__a22o_2 _09805_ (.A1(_03698_),
    .A2(_04059_),
    .B1(_04060_),
    .B2(_03686_),
    .X(_04061_));
 sky130_fd_sc_hd__o211a_2 _09806_ (.A1(_03679_),
    .A2(\core.reg_next_pc[31] ),
    .B1(_03915_),
    .C1(_04061_),
    .X(_00147_));
 sky130_fd_sc_hd__a22o_2 _09807_ (.A1(_03713_),
    .A2(_03658_),
    .B1(_03780_),
    .B2(\core.reg_pc[1] ),
    .X(_00148_));
 sky130_fd_sc_hd__a22o_2 _09808_ (.A1(_03713_),
    .A2(_03670_),
    .B1(_03780_),
    .B2(_02493_),
    .X(_00149_));
 sky130_fd_sc_hd__o211a_2 _09809_ (.A1(_03679_),
    .A2(\core.reg_pc[3] ),
    .B1(_03915_),
    .C1(_03684_),
    .X(_00150_));
 sky130_fd_sc_hd__buf_1 _09810_ (.A(_02080_),
    .X(_04062_));
 sky130_fd_sc_hd__o211a_2 _09811_ (.A1(_04062_),
    .A2(\core.reg_pc[4] ),
    .B1(_03915_),
    .C1(_03711_),
    .X(_00151_));
 sky130_fd_sc_hd__buf_1 _09812_ (.A(_02111_),
    .X(_04063_));
 sky130_fd_sc_hd__a22o_2 _09813_ (.A1(\core.reg_pc[5] ),
    .A2(_03780_),
    .B1(_03717_),
    .B2(_04063_),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_2 _09814_ (.A1(\core.reg_pc[6] ),
    .A2(_03780_),
    .B1(_03731_),
    .B2(_04063_),
    .X(_00153_));
 sky130_fd_sc_hd__o211a_2 _09815_ (.A1(_04062_),
    .A2(\core.reg_pc[7] ),
    .B1(_03915_),
    .C1(_03748_),
    .X(_00154_));
 sky130_fd_sc_hd__o211a_2 _09816_ (.A1(_04062_),
    .A2(\core.reg_pc[8] ),
    .B1(_03915_),
    .C1(_03762_),
    .X(_00155_));
 sky130_fd_sc_hd__a22o_2 _09817_ (.A1(\core.reg_pc[9] ),
    .A2(_03780_),
    .B1(_03771_),
    .B2(_04063_),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_2 _09818_ (.A1(\core.reg_pc[10] ),
    .A2(_03780_),
    .B1(_03782_),
    .B2(_04063_),
    .X(_00157_));
 sky130_fd_sc_hd__o211a_2 _09819_ (.A1(_04062_),
    .A2(\core.reg_pc[11] ),
    .B1(_03915_),
    .C1(_03804_),
    .X(_00158_));
 sky130_fd_sc_hd__o211a_2 _09820_ (.A1(_04062_),
    .A2(\core.reg_pc[12] ),
    .B1(_03915_),
    .C1(_03817_),
    .X(_00159_));
 sky130_fd_sc_hd__a22o_2 _09821_ (.A1(\core.reg_pc[13] ),
    .A2(_03780_),
    .B1(_03827_),
    .B2(_04063_),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_2 _09822_ (.A1(\core.reg_pc[14] ),
    .A2(_03780_),
    .B1(_03837_),
    .B2(_04063_),
    .X(_00161_));
 sky130_fd_sc_hd__o211a_2 _09823_ (.A1(_04062_),
    .A2(\core.reg_pc[15] ),
    .B1(_02083_),
    .C1(_03856_),
    .X(_00162_));
 sky130_fd_sc_hd__or2_2 _09824_ (.A(_02080_),
    .B(\core.reg_pc[16] ),
    .X(_04064_));
 sky130_fd_sc_hd__o211a_2 _09825_ (.A1(_03663_),
    .A2(_03864_),
    .B1(_04064_),
    .C1(_03665_),
    .X(_00163_));
 sky130_fd_sc_hd__a22o_2 _09826_ (.A1(\core.reg_pc[17] ),
    .A2(_03729_),
    .B1(_03882_),
    .B2(_04063_),
    .X(_00164_));
 sky130_fd_sc_hd__a22o_2 _09827_ (.A1(\core.reg_pc[18] ),
    .A2(_03729_),
    .B1(_03893_),
    .B2(_04063_),
    .X(_00165_));
 sky130_fd_sc_hd__o211a_2 _09828_ (.A1(_04062_),
    .A2(\core.reg_pc[19] ),
    .B1(_02083_),
    .C1(_03910_),
    .X(_00166_));
 sky130_fd_sc_hd__o211a_2 _09829_ (.A1(_04062_),
    .A2(\core.reg_pc[20] ),
    .B1(_02083_),
    .C1(_03926_),
    .X(_00167_));
 sky130_fd_sc_hd__a22o_2 _09830_ (.A1(\core.reg_pc[21] ),
    .A2(_03729_),
    .B1(_03929_),
    .B2(_04063_),
    .X(_00168_));
 sky130_fd_sc_hd__or2_2 _09831_ (.A(_02080_),
    .B(\core.reg_pc[22] ),
    .X(_04065_));
 sky130_fd_sc_hd__o211a_2 _09832_ (.A1(_03663_),
    .A2(_03946_),
    .B1(_04065_),
    .C1(_03665_),
    .X(_00169_));
 sky130_fd_sc_hd__o211a_2 _09833_ (.A1(_04062_),
    .A2(\core.reg_pc[23] ),
    .B1(_02083_),
    .C1(_03958_),
    .X(_00170_));
 sky130_fd_sc_hd__or2_2 _09834_ (.A(_02080_),
    .B(\core.reg_pc[24] ),
    .X(_04066_));
 sky130_fd_sc_hd__o211a_2 _09835_ (.A1(_03663_),
    .A2(_03972_),
    .B1(_04066_),
    .C1(_03665_),
    .X(_00171_));
 sky130_fd_sc_hd__a22o_2 _09836_ (.A1(\core.reg_pc[25] ),
    .A2(_03729_),
    .B1(_03989_),
    .B2(_04063_),
    .X(_00172_));
 sky130_fd_sc_hd__o211a_2 _09837_ (.A1(_04062_),
    .A2(\core.reg_pc[26] ),
    .B1(_02083_),
    .C1(_04006_),
    .X(_00173_));
 sky130_fd_sc_hd__a22o_2 _09838_ (.A1(\core.reg_pc[27] ),
    .A2(_03729_),
    .B1(_04011_),
    .B2(_03713_),
    .X(_00174_));
 sky130_fd_sc_hd__o211a_2 _09839_ (.A1(_03655_),
    .A2(\core.reg_pc[28] ),
    .B1(_02083_),
    .C1(_04027_),
    .X(_00175_));
 sky130_fd_sc_hd__a22o_2 _09840_ (.A1(\core.reg_pc[29] ),
    .A2(_03729_),
    .B1(_04032_),
    .B2(_03713_),
    .X(_00176_));
 sky130_fd_sc_hd__o211a_2 _09841_ (.A1(_03655_),
    .A2(\core.reg_pc[30] ),
    .B1(_02083_),
    .C1(_04051_),
    .X(_00177_));
 sky130_fd_sc_hd__o211a_2 _09842_ (.A1(\core.reg_pc[31] ),
    .A2(_03679_),
    .B1(_02083_),
    .C1(_04060_),
    .X(_00178_));
 sky130_fd_sc_hd__and3_2 _09843_ (.A(\core.count_instr[0] ),
    .B(_02079_),
    .C(_03659_),
    .X(_04067_));
 sky130_fd_sc_hd__a21o_2 _09844_ (.A1(_02079_),
    .A2(_03659_),
    .B1(\core.count_instr[0] ),
    .X(_04068_));
 sky130_fd_sc_hd__and3b_2 _09845_ (.A_N(_04067_),
    .B(_04068_),
    .C(_02082_),
    .X(_04069_));
 sky130_fd_sc_hd__buf_1 _09846_ (.A(_04069_),
    .X(_00179_));
 sky130_fd_sc_hd__and4_2 _09847_ (.A(\core.count_instr[1] ),
    .B(\core.count_instr[0] ),
    .C(\core.cpu_state[1] ),
    .D(\core.decoder_trigger ),
    .X(_04070_));
 sky130_fd_sc_hd__o21ai_2 _09848_ (.A1(\core.count_instr[1] ),
    .A2(_04067_),
    .B1(_03482_),
    .Y(_04071_));
 sky130_fd_sc_hd__nor2_2 _09849_ (.A(_04070_),
    .B(_04071_),
    .Y(_00180_));
 sky130_fd_sc_hd__a21oi_2 _09850_ (.A1(\core.count_instr[2] ),
    .A2(_04070_),
    .B1(_03498_),
    .Y(_04072_));
 sky130_fd_sc_hd__o21a_2 _09851_ (.A1(\core.count_instr[2] ),
    .A2(_04070_),
    .B1(_04072_),
    .X(_00181_));
 sky130_fd_sc_hd__and3_2 _09852_ (.A(\core.count_instr[3] ),
    .B(\core.count_instr[2] ),
    .C(_04070_),
    .X(_04073_));
 sky130_fd_sc_hd__a21o_2 _09853_ (.A1(\core.count_instr[2] ),
    .A2(_04070_),
    .B1(\core.count_instr[3] ),
    .X(_04074_));
 sky130_fd_sc_hd__and3b_2 _09854_ (.A_N(_04073_),
    .B(_03621_),
    .C(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__buf_1 _09855_ (.A(_04075_),
    .X(_00182_));
 sky130_fd_sc_hd__o21ai_2 _09856_ (.A1(\core.count_instr[4] ),
    .A2(_04073_),
    .B1(_03482_),
    .Y(_04076_));
 sky130_fd_sc_hd__a21oi_2 _09857_ (.A1(\core.count_instr[4] ),
    .A2(_04073_),
    .B1(_04076_),
    .Y(_00183_));
 sky130_fd_sc_hd__and2_2 _09858_ (.A(\core.count_instr[5] ),
    .B(\core.count_instr[4] ),
    .X(_04077_));
 sky130_fd_sc_hd__and4_2 _09859_ (.A(\core.count_instr[3] ),
    .B(\core.count_instr[2] ),
    .C(_04070_),
    .D(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__a21o_2 _09860_ (.A1(\core.count_instr[4] ),
    .A2(_04073_),
    .B1(\core.count_instr[5] ),
    .X(_04079_));
 sky130_fd_sc_hd__and3b_2 _09861_ (.A_N(_04078_),
    .B(_03621_),
    .C(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__buf_1 _09862_ (.A(_04080_),
    .X(_00184_));
 sky130_fd_sc_hd__and2_2 _09863_ (.A(\core.count_instr[6] ),
    .B(_04078_),
    .X(_04081_));
 sky130_fd_sc_hd__nor2_2 _09864_ (.A(_03557_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__o21a_2 _09865_ (.A1(\core.count_instr[6] ),
    .A2(_04078_),
    .B1(_04082_),
    .X(_00185_));
 sky130_fd_sc_hd__and3_2 _09866_ (.A(\core.count_instr[7] ),
    .B(\core.count_instr[6] ),
    .C(_04078_),
    .X(_04083_));
 sky130_fd_sc_hd__or2_2 _09867_ (.A(\core.count_instr[7] ),
    .B(_04081_),
    .X(_04084_));
 sky130_fd_sc_hd__and3b_2 _09868_ (.A_N(_04083_),
    .B(_03621_),
    .C(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__buf_1 _09869_ (.A(_04085_),
    .X(_00186_));
 sky130_fd_sc_hd__o21ai_2 _09870_ (.A1(\core.count_instr[8] ),
    .A2(_04083_),
    .B1(_03482_),
    .Y(_04086_));
 sky130_fd_sc_hd__a21oi_2 _09871_ (.A1(\core.count_instr[8] ),
    .A2(_04083_),
    .B1(_04086_),
    .Y(_00187_));
 sky130_fd_sc_hd__and2_2 _09872_ (.A(\core.count_instr[9] ),
    .B(\core.count_instr[8] ),
    .X(_04087_));
 sky130_fd_sc_hd__and4_2 _09873_ (.A(\core.count_instr[7] ),
    .B(\core.count_instr[6] ),
    .C(_04078_),
    .D(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__a21o_2 _09874_ (.A1(\core.count_instr[8] ),
    .A2(_04083_),
    .B1(\core.count_instr[9] ),
    .X(_04089_));
 sky130_fd_sc_hd__and3b_2 _09875_ (.A_N(_04088_),
    .B(_03621_),
    .C(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__buf_1 _09876_ (.A(_04090_),
    .X(_00188_));
 sky130_fd_sc_hd__and2_2 _09877_ (.A(\core.count_instr[10] ),
    .B(_04088_),
    .X(_04091_));
 sky130_fd_sc_hd__nor2_2 _09878_ (.A(_03557_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__o21a_2 _09879_ (.A1(\core.count_instr[10] ),
    .A2(_04088_),
    .B1(_04092_),
    .X(_00189_));
 sky130_fd_sc_hd__and3_2 _09880_ (.A(\core.count_instr[11] ),
    .B(\core.count_instr[10] ),
    .C(_04088_),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_2 _09881_ (.A(_03557_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__o21a_2 _09882_ (.A1(\core.count_instr[11] ),
    .A2(_04091_),
    .B1(_04094_),
    .X(_00190_));
 sky130_fd_sc_hd__o21ai_2 _09883_ (.A1(\core.count_instr[12] ),
    .A2(_04093_),
    .B1(_03482_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_2 _09884_ (.A1(\core.count_instr[12] ),
    .A2(_04093_),
    .B1(_04095_),
    .Y(_00191_));
 sky130_fd_sc_hd__and2_2 _09885_ (.A(\core.count_instr[13] ),
    .B(\core.count_instr[12] ),
    .X(_04096_));
 sky130_fd_sc_hd__and4_2 _09886_ (.A(\core.count_instr[11] ),
    .B(\core.count_instr[10] ),
    .C(_04088_),
    .D(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__a21o_2 _09887_ (.A1(\core.count_instr[12] ),
    .A2(_04093_),
    .B1(\core.count_instr[13] ),
    .X(_04098_));
 sky130_fd_sc_hd__and3b_2 _09888_ (.A_N(_04097_),
    .B(_03621_),
    .C(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__buf_1 _09889_ (.A(_04099_),
    .X(_00192_));
 sky130_fd_sc_hd__and2_2 _09890_ (.A(\core.count_instr[14] ),
    .B(_04097_),
    .X(_04100_));
 sky130_fd_sc_hd__nor2_2 _09891_ (.A(_03557_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__o21a_2 _09892_ (.A1(\core.count_instr[14] ),
    .A2(_04097_),
    .B1(_04101_),
    .X(_00193_));
 sky130_fd_sc_hd__and3_2 _09893_ (.A(\core.count_instr[15] ),
    .B(\core.count_instr[14] ),
    .C(_04097_),
    .X(_04102_));
 sky130_fd_sc_hd__buf_1 _09894_ (.A(_02024_),
    .X(_04103_));
 sky130_fd_sc_hd__or2_2 _09895_ (.A(\core.count_instr[15] ),
    .B(_04100_),
    .X(_04104_));
 sky130_fd_sc_hd__and3b_2 _09896_ (.A_N(_04102_),
    .B(_04103_),
    .C(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__buf_1 _09897_ (.A(_04105_),
    .X(_00194_));
 sky130_fd_sc_hd__o21ai_2 _09898_ (.A1(\core.count_instr[16] ),
    .A2(_04102_),
    .B1(_03482_),
    .Y(_04106_));
 sky130_fd_sc_hd__a21oi_2 _09899_ (.A1(\core.count_instr[16] ),
    .A2(_04102_),
    .B1(_04106_),
    .Y(_00195_));
 sky130_fd_sc_hd__and2_2 _09900_ (.A(\core.count_instr[17] ),
    .B(\core.count_instr[16] ),
    .X(_04107_));
 sky130_fd_sc_hd__and4_2 _09901_ (.A(\core.count_instr[15] ),
    .B(\core.count_instr[14] ),
    .C(_04097_),
    .D(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__a21o_2 _09902_ (.A1(\core.count_instr[16] ),
    .A2(_04102_),
    .B1(\core.count_instr[17] ),
    .X(_04109_));
 sky130_fd_sc_hd__and3b_2 _09903_ (.A_N(_04108_),
    .B(_04103_),
    .C(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__buf_1 _09904_ (.A(_04110_),
    .X(_00196_));
 sky130_fd_sc_hd__and2_2 _09905_ (.A(\core.count_instr[18] ),
    .B(_04108_),
    .X(_04111_));
 sky130_fd_sc_hd__nor2_2 _09906_ (.A(_03557_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__o21a_2 _09907_ (.A1(\core.count_instr[18] ),
    .A2(_04108_),
    .B1(_04112_),
    .X(_00197_));
 sky130_fd_sc_hd__and3_2 _09908_ (.A(\core.count_instr[19] ),
    .B(\core.count_instr[18] ),
    .C(_04108_),
    .X(_04113_));
 sky130_fd_sc_hd__or2_2 _09909_ (.A(\core.count_instr[19] ),
    .B(_04111_),
    .X(_04114_));
 sky130_fd_sc_hd__and3b_2 _09910_ (.A_N(_04113_),
    .B(_04103_),
    .C(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__buf_1 _09911_ (.A(_04115_),
    .X(_00198_));
 sky130_fd_sc_hd__o21ai_2 _09912_ (.A1(\core.count_instr[20] ),
    .A2(_04113_),
    .B1(_03482_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21oi_2 _09913_ (.A1(\core.count_instr[20] ),
    .A2(_04113_),
    .B1(_04116_),
    .Y(_00199_));
 sky130_fd_sc_hd__and2_2 _09914_ (.A(\core.count_instr[21] ),
    .B(\core.count_instr[20] ),
    .X(_04117_));
 sky130_fd_sc_hd__and4_2 _09915_ (.A(\core.count_instr[19] ),
    .B(\core.count_instr[18] ),
    .C(_04108_),
    .D(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__a21o_2 _09916_ (.A1(\core.count_instr[20] ),
    .A2(_04113_),
    .B1(\core.count_instr[21] ),
    .X(_04119_));
 sky130_fd_sc_hd__and3b_2 _09917_ (.A_N(_04118_),
    .B(_04103_),
    .C(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__buf_1 _09918_ (.A(_04120_),
    .X(_00200_));
 sky130_fd_sc_hd__buf_1 _09919_ (.A(_02049_),
    .X(_04121_));
 sky130_fd_sc_hd__and2_2 _09920_ (.A(\core.count_instr[22] ),
    .B(_04118_),
    .X(_04122_));
 sky130_fd_sc_hd__nor2_2 _09921_ (.A(_04121_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__o21a_2 _09922_ (.A1(\core.count_instr[22] ),
    .A2(_04118_),
    .B1(_04123_),
    .X(_00201_));
 sky130_fd_sc_hd__and3_2 _09923_ (.A(\core.count_instr[23] ),
    .B(\core.count_instr[22] ),
    .C(_04118_),
    .X(_04124_));
 sky130_fd_sc_hd__nor2_2 _09924_ (.A(_04121_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__o21a_2 _09925_ (.A1(\core.count_instr[23] ),
    .A2(_04122_),
    .B1(_04125_),
    .X(_00202_));
 sky130_fd_sc_hd__o21ai_2 _09926_ (.A1(\core.count_instr[24] ),
    .A2(_04124_),
    .B1(_03482_),
    .Y(_04126_));
 sky130_fd_sc_hd__a21oi_2 _09927_ (.A1(\core.count_instr[24] ),
    .A2(_04124_),
    .B1(_04126_),
    .Y(_00203_));
 sky130_fd_sc_hd__and2_2 _09928_ (.A(\core.count_instr[25] ),
    .B(\core.count_instr[24] ),
    .X(_04127_));
 sky130_fd_sc_hd__and4_2 _09929_ (.A(\core.count_instr[23] ),
    .B(\core.count_instr[22] ),
    .C(_04118_),
    .D(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__a21o_2 _09930_ (.A1(\core.count_instr[24] ),
    .A2(_04124_),
    .B1(\core.count_instr[25] ),
    .X(_04129_));
 sky130_fd_sc_hd__and3b_2 _09931_ (.A_N(_04128_),
    .B(_04103_),
    .C(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__buf_1 _09932_ (.A(_04130_),
    .X(_00204_));
 sky130_fd_sc_hd__and2_2 _09933_ (.A(\core.count_instr[26] ),
    .B(_04128_),
    .X(_04131_));
 sky130_fd_sc_hd__nor2_2 _09934_ (.A(_04121_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__o21a_2 _09935_ (.A1(\core.count_instr[26] ),
    .A2(_04128_),
    .B1(_04132_),
    .X(_00205_));
 sky130_fd_sc_hd__and3_2 _09936_ (.A(\core.count_instr[27] ),
    .B(\core.count_instr[26] ),
    .C(_04128_),
    .X(_04133_));
 sky130_fd_sc_hd__nor2_2 _09937_ (.A(_04121_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21a_2 _09938_ (.A1(\core.count_instr[27] ),
    .A2(_04131_),
    .B1(_04134_),
    .X(_00206_));
 sky130_fd_sc_hd__o21ai_2 _09939_ (.A1(\core.count_instr[28] ),
    .A2(_04133_),
    .B1(_03482_),
    .Y(_04135_));
 sky130_fd_sc_hd__a21oi_2 _09940_ (.A1(\core.count_instr[28] ),
    .A2(_04133_),
    .B1(_04135_),
    .Y(_00207_));
 sky130_fd_sc_hd__and2_2 _09941_ (.A(\core.count_instr[29] ),
    .B(\core.count_instr[28] ),
    .X(_04136_));
 sky130_fd_sc_hd__and4_2 _09942_ (.A(\core.count_instr[27] ),
    .B(\core.count_instr[26] ),
    .C(_04128_),
    .D(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__a21o_2 _09943_ (.A1(\core.count_instr[28] ),
    .A2(_04133_),
    .B1(\core.count_instr[29] ),
    .X(_04138_));
 sky130_fd_sc_hd__and3b_2 _09944_ (.A_N(_04137_),
    .B(_04103_),
    .C(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__buf_1 _09945_ (.A(_04139_),
    .X(_00208_));
 sky130_fd_sc_hd__and2_2 _09946_ (.A(\core.count_instr[30] ),
    .B(_04137_),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_2 _09947_ (.A(_04121_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__o21a_2 _09948_ (.A1(\core.count_instr[30] ),
    .A2(_04137_),
    .B1(_04141_),
    .X(_00209_));
 sky130_fd_sc_hd__and3_2 _09949_ (.A(\core.count_instr[31] ),
    .B(\core.count_instr[30] ),
    .C(_04137_),
    .X(_04142_));
 sky130_fd_sc_hd__nor2_2 _09950_ (.A(_04121_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__o21a_2 _09951_ (.A1(\core.count_instr[31] ),
    .A2(_04140_),
    .B1(_04143_),
    .X(_00210_));
 sky130_fd_sc_hd__buf_1 _09952_ (.A(_02052_),
    .X(_04144_));
 sky130_fd_sc_hd__o21ai_2 _09953_ (.A1(\core.count_instr[32] ),
    .A2(_04142_),
    .B1(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a21oi_2 _09954_ (.A1(\core.count_instr[32] ),
    .A2(_04142_),
    .B1(_04145_),
    .Y(_00211_));
 sky130_fd_sc_hd__and2_2 _09955_ (.A(\core.count_instr[33] ),
    .B(\core.count_instr[32] ),
    .X(_04146_));
 sky130_fd_sc_hd__and4_2 _09956_ (.A(\core.count_instr[31] ),
    .B(\core.count_instr[30] ),
    .C(_04137_),
    .D(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__a21o_2 _09957_ (.A1(\core.count_instr[32] ),
    .A2(_04142_),
    .B1(\core.count_instr[33] ),
    .X(_04148_));
 sky130_fd_sc_hd__and3b_2 _09958_ (.A_N(_04147_),
    .B(_04103_),
    .C(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__buf_1 _09959_ (.A(_04149_),
    .X(_00212_));
 sky130_fd_sc_hd__and2_2 _09960_ (.A(\core.count_instr[34] ),
    .B(_04147_),
    .X(_04150_));
 sky130_fd_sc_hd__nor2_2 _09961_ (.A(_04121_),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__o21a_2 _09962_ (.A1(\core.count_instr[34] ),
    .A2(_04147_),
    .B1(_04151_),
    .X(_00213_));
 sky130_fd_sc_hd__and3_2 _09963_ (.A(\core.count_instr[35] ),
    .B(\core.count_instr[34] ),
    .C(_04147_),
    .X(_04152_));
 sky130_fd_sc_hd__nor2_2 _09964_ (.A(_04121_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__o21a_2 _09965_ (.A1(\core.count_instr[35] ),
    .A2(_04150_),
    .B1(_04153_),
    .X(_00214_));
 sky130_fd_sc_hd__o21ai_2 _09966_ (.A1(\core.count_instr[36] ),
    .A2(_04152_),
    .B1(_04144_),
    .Y(_04154_));
 sky130_fd_sc_hd__a21oi_2 _09967_ (.A1(\core.count_instr[36] ),
    .A2(_04152_),
    .B1(_04154_),
    .Y(_00215_));
 sky130_fd_sc_hd__and2_2 _09968_ (.A(\core.count_instr[37] ),
    .B(\core.count_instr[36] ),
    .X(_04155_));
 sky130_fd_sc_hd__and4_2 _09969_ (.A(\core.count_instr[35] ),
    .B(\core.count_instr[34] ),
    .C(_04147_),
    .D(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__a21o_2 _09970_ (.A1(\core.count_instr[36] ),
    .A2(_04152_),
    .B1(\core.count_instr[37] ),
    .X(_04157_));
 sky130_fd_sc_hd__and3b_2 _09971_ (.A_N(_04156_),
    .B(_04103_),
    .C(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__buf_1 _09972_ (.A(_04158_),
    .X(_00216_));
 sky130_fd_sc_hd__and2_2 _09973_ (.A(\core.count_instr[38] ),
    .B(_04156_),
    .X(_04159_));
 sky130_fd_sc_hd__nor2_2 _09974_ (.A(_04121_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__o21a_2 _09975_ (.A1(\core.count_instr[38] ),
    .A2(_04156_),
    .B1(_04160_),
    .X(_00217_));
 sky130_fd_sc_hd__and3_2 _09976_ (.A(\core.count_instr[39] ),
    .B(\core.count_instr[38] ),
    .C(_04156_),
    .X(_04161_));
 sky130_fd_sc_hd__nor2_2 _09977_ (.A(_04121_),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__o21a_2 _09978_ (.A1(\core.count_instr[39] ),
    .A2(_04159_),
    .B1(_04162_),
    .X(_00218_));
 sky130_fd_sc_hd__o21ai_2 _09979_ (.A1(\core.count_instr[40] ),
    .A2(_04161_),
    .B1(_04144_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_2 _09980_ (.A1(\core.count_instr[40] ),
    .A2(_04161_),
    .B1(_04163_),
    .Y(_00219_));
 sky130_fd_sc_hd__and2_2 _09981_ (.A(\core.count_instr[41] ),
    .B(\core.count_instr[40] ),
    .X(_04164_));
 sky130_fd_sc_hd__and4_2 _09982_ (.A(\core.count_instr[39] ),
    .B(\core.count_instr[38] ),
    .C(_04156_),
    .D(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__a21o_2 _09983_ (.A1(\core.count_instr[40] ),
    .A2(_04161_),
    .B1(\core.count_instr[41] ),
    .X(_04166_));
 sky130_fd_sc_hd__and3b_2 _09984_ (.A_N(_04165_),
    .B(_04103_),
    .C(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__buf_1 _09985_ (.A(_04167_),
    .X(_00220_));
 sky130_fd_sc_hd__nand2_2 _09986_ (.A(\core.count_instr[42] ),
    .B(_04165_),
    .Y(_04168_));
 sky130_fd_sc_hd__and2_2 _09987_ (.A(_02082_),
    .B(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__o21a_2 _09988_ (.A1(\core.count_instr[42] ),
    .A2(_04165_),
    .B1(_04169_),
    .X(_00221_));
 sky130_fd_sc_hd__inv_2 _09989_ (.A(\core.count_instr[43] ),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_2 _09990_ (.A(_04170_),
    .B(_04168_),
    .Y(_04171_));
 sky130_fd_sc_hd__or2_2 _09991_ (.A(_02049_),
    .B(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__a21oi_2 _09992_ (.A1(_04170_),
    .A2(_04168_),
    .B1(_04172_),
    .Y(_00222_));
 sky130_fd_sc_hd__o21ai_2 _09993_ (.A1(\core.count_instr[44] ),
    .A2(_04171_),
    .B1(_04144_),
    .Y(_04173_));
 sky130_fd_sc_hd__a21oi_2 _09994_ (.A1(\core.count_instr[44] ),
    .A2(_04171_),
    .B1(_04173_),
    .Y(_00223_));
 sky130_fd_sc_hd__and2_2 _09995_ (.A(\core.count_instr[45] ),
    .B(\core.count_instr[44] ),
    .X(_04174_));
 sky130_fd_sc_hd__and4_2 _09996_ (.A(\core.count_instr[43] ),
    .B(\core.count_instr[42] ),
    .C(_04165_),
    .D(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__a21o_2 _09997_ (.A1(\core.count_instr[44] ),
    .A2(_04171_),
    .B1(\core.count_instr[45] ),
    .X(_04176_));
 sky130_fd_sc_hd__and3b_2 _09998_ (.A_N(_04175_),
    .B(_04103_),
    .C(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__buf_1 _09999_ (.A(_04177_),
    .X(_00224_));
 sky130_fd_sc_hd__and2_2 _10000_ (.A(\core.count_instr[46] ),
    .B(_04175_),
    .X(_04178_));
 sky130_fd_sc_hd__nor2_2 _10001_ (.A(_02054_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__o21a_2 _10002_ (.A1(\core.count_instr[46] ),
    .A2(_04175_),
    .B1(_04179_),
    .X(_00225_));
 sky130_fd_sc_hd__and3_2 _10003_ (.A(\core.count_instr[47] ),
    .B(\core.count_instr[46] ),
    .C(_04175_),
    .X(_04180_));
 sky130_fd_sc_hd__nor2_2 _10004_ (.A(_02054_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__o21a_2 _10005_ (.A1(\core.count_instr[47] ),
    .A2(_04178_),
    .B1(_04181_),
    .X(_00226_));
 sky130_fd_sc_hd__o21ai_2 _10006_ (.A1(\core.count_instr[48] ),
    .A2(_04180_),
    .B1(_04144_),
    .Y(_04182_));
 sky130_fd_sc_hd__a21oi_2 _10007_ (.A1(\core.count_instr[48] ),
    .A2(_04180_),
    .B1(_04182_),
    .Y(_00227_));
 sky130_fd_sc_hd__and2_2 _10008_ (.A(\core.count_instr[49] ),
    .B(\core.count_instr[48] ),
    .X(_04183_));
 sky130_fd_sc_hd__and4_2 _10009_ (.A(\core.count_instr[47] ),
    .B(\core.count_instr[46] ),
    .C(_04175_),
    .D(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__a21o_2 _10010_ (.A1(\core.count_instr[48] ),
    .A2(_04180_),
    .B1(\core.count_instr[49] ),
    .X(_04185_));
 sky130_fd_sc_hd__and3b_2 _10011_ (.A_N(_04184_),
    .B(_02082_),
    .C(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__buf_1 _10012_ (.A(_04186_),
    .X(_00228_));
 sky130_fd_sc_hd__and2_2 _10013_ (.A(\core.count_instr[50] ),
    .B(_04184_),
    .X(_04187_));
 sky130_fd_sc_hd__nor2_2 _10014_ (.A(_02054_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__o21a_2 _10015_ (.A1(\core.count_instr[50] ),
    .A2(_04184_),
    .B1(_04188_),
    .X(_00229_));
 sky130_fd_sc_hd__and3_2 _10016_ (.A(\core.count_instr[51] ),
    .B(\core.count_instr[50] ),
    .C(_04184_),
    .X(_04189_));
 sky130_fd_sc_hd__nor2_2 _10017_ (.A(_02054_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__o21a_2 _10018_ (.A1(\core.count_instr[51] ),
    .A2(_04187_),
    .B1(_04190_),
    .X(_00230_));
 sky130_fd_sc_hd__and4_2 _10019_ (.A(\core.count_instr[52] ),
    .B(\core.count_instr[51] ),
    .C(\core.count_instr[50] ),
    .D(_04184_),
    .X(_04191_));
 sky130_fd_sc_hd__nor2_2 _10020_ (.A(_02054_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__o21a_2 _10021_ (.A1(\core.count_instr[52] ),
    .A2(_04189_),
    .B1(_04192_),
    .X(_00231_));
 sky130_fd_sc_hd__or2_2 _10022_ (.A(\core.count_instr[53] ),
    .B(_04191_),
    .X(_04193_));
 sky130_fd_sc_hd__nand2_2 _10023_ (.A(\core.count_instr[53] ),
    .B(_04191_),
    .Y(_04194_));
 sky130_fd_sc_hd__and3_2 _10024_ (.A(_03571_),
    .B(_04193_),
    .C(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__buf_1 _10025_ (.A(_04195_),
    .X(_00232_));
 sky130_fd_sc_hd__inv_2 _10026_ (.A(\core.count_instr[54] ),
    .Y(_04196_));
 sky130_fd_sc_hd__a31o_2 _10027_ (.A1(\core.count_instr[54] ),
    .A2(\core.count_instr[53] ),
    .A3(_04191_),
    .B1(_02049_),
    .X(_04197_));
 sky130_fd_sc_hd__a21oi_2 _10028_ (.A1(_04196_),
    .A2(_04194_),
    .B1(_04197_),
    .Y(_00233_));
 sky130_fd_sc_hd__and4_2 _10029_ (.A(\core.count_instr[55] ),
    .B(\core.count_instr[54] ),
    .C(\core.count_instr[53] ),
    .D(_04191_),
    .X(_04198_));
 sky130_fd_sc_hd__a31o_2 _10030_ (.A1(\core.count_instr[54] ),
    .A2(\core.count_instr[53] ),
    .A3(_04191_),
    .B1(\core.count_instr[55] ),
    .X(_04199_));
 sky130_fd_sc_hd__and3b_2 _10031_ (.A_N(_04198_),
    .B(_02082_),
    .C(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__buf_1 _10032_ (.A(_04200_),
    .X(_00234_));
 sky130_fd_sc_hd__a21oi_2 _10033_ (.A1(\core.count_instr[56] ),
    .A2(_04198_),
    .B1(_03498_),
    .Y(_04201_));
 sky130_fd_sc_hd__o21a_2 _10034_ (.A1(\core.count_instr[56] ),
    .A2(_04198_),
    .B1(_04201_),
    .X(_00235_));
 sky130_fd_sc_hd__and3_2 _10035_ (.A(\core.count_instr[57] ),
    .B(\core.count_instr[56] ),
    .C(_04198_),
    .X(_04202_));
 sky130_fd_sc_hd__a21o_2 _10036_ (.A1(\core.count_instr[56] ),
    .A2(_04198_),
    .B1(\core.count_instr[57] ),
    .X(_04203_));
 sky130_fd_sc_hd__and3b_2 _10037_ (.A_N(_04202_),
    .B(_02082_),
    .C(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__buf_1 _10038_ (.A(_04204_),
    .X(_00236_));
 sky130_fd_sc_hd__and4_2 _10039_ (.A(\core.count_instr[58] ),
    .B(\core.count_instr[57] ),
    .C(\core.count_instr[56] ),
    .D(_04198_),
    .X(_04205_));
 sky130_fd_sc_hd__nor2_2 _10040_ (.A(_02054_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__o21a_2 _10041_ (.A1(\core.count_instr[58] ),
    .A2(_04202_),
    .B1(_04206_),
    .X(_00237_));
 sky130_fd_sc_hd__a21oi_2 _10042_ (.A1(\core.count_instr[59] ),
    .A2(_04205_),
    .B1(_03498_),
    .Y(_04207_));
 sky130_fd_sc_hd__o21a_2 _10043_ (.A1(\core.count_instr[59] ),
    .A2(_04205_),
    .B1(_04207_),
    .X(_00238_));
 sky130_fd_sc_hd__and3_2 _10044_ (.A(\core.count_instr[60] ),
    .B(\core.count_instr[59] ),
    .C(_04205_),
    .X(_04208_));
 sky130_fd_sc_hd__a21o_2 _10045_ (.A1(\core.count_instr[59] ),
    .A2(_04205_),
    .B1(\core.count_instr[60] ),
    .X(_04209_));
 sky130_fd_sc_hd__and3b_2 _10046_ (.A_N(_04208_),
    .B(_02082_),
    .C(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__buf_1 _10047_ (.A(_04210_),
    .X(_00239_));
 sky130_fd_sc_hd__and4_2 _10048_ (.A(\core.count_instr[61] ),
    .B(\core.count_instr[60] ),
    .C(\core.count_instr[59] ),
    .D(_04205_),
    .X(_04211_));
 sky130_fd_sc_hd__nor2_2 _10049_ (.A(_02054_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__o21a_2 _10050_ (.A1(\core.count_instr[61] ),
    .A2(_04208_),
    .B1(_04212_),
    .X(_00240_));
 sky130_fd_sc_hd__a21oi_2 _10051_ (.A1(\core.count_instr[62] ),
    .A2(_04211_),
    .B1(_03498_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21a_2 _10052_ (.A1(\core.count_instr[62] ),
    .A2(_04211_),
    .B1(_04213_),
    .X(_00241_));
 sky130_fd_sc_hd__nand3_2 _10053_ (.A(\core.count_instr[63] ),
    .B(\core.count_instr[62] ),
    .C(_04211_),
    .Y(_04214_));
 sky130_fd_sc_hd__a21o_2 _10054_ (.A1(\core.count_instr[62] ),
    .A2(_04211_),
    .B1(\core.count_instr[63] ),
    .X(_04215_));
 sky130_fd_sc_hd__and3_2 _10055_ (.A(_03571_),
    .B(_04214_),
    .C(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_1 _10056_ (.A(_04216_),
    .X(_00242_));
 sky130_fd_sc_hd__buf_1 _10057_ (.A(_03271_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_1 _10058_ (.A(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__buf_1 _10059_ (.A(_03277_),
    .X(_04219_));
 sky130_fd_sc_hd__buf_1 _10060_ (.A(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__mux4_2 _10061_ (.A0(\core.cpuregs[20][0] ),
    .A1(\core.cpuregs[21][0] ),
    .A2(\core.cpuregs[22][0] ),
    .A3(\core.cpuregs[23][0] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__mux4_2 _10062_ (.A0(\core.cpuregs[16][0] ),
    .A1(\core.cpuregs[17][0] ),
    .A2(\core.cpuregs[18][0] ),
    .A3(\core.cpuregs[19][0] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_04222_));
 sky130_fd_sc_hd__mux2_2 _10063_ (.A0(_04221_),
    .A1(_04222_),
    .S(_03295_),
    .X(_04223_));
 sky130_fd_sc_hd__buf_1 _10064_ (.A(_04219_),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_2 _10065_ (.A0(\core.cpuregs[28][0] ),
    .A1(\core.cpuregs[29][0] ),
    .A2(\core.cpuregs[30][0] ),
    .A3(\core.cpuregs[31][0] ),
    .S0(_04218_),
    .S1(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__mux4_2 _10066_ (.A0(\core.cpuregs[24][0] ),
    .A1(\core.cpuregs[25][0] ),
    .A2(\core.cpuregs[26][0] ),
    .A3(\core.cpuregs[27][0] ),
    .S0(_04218_),
    .S1(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__mux2_2 _10067_ (.A0(_04225_),
    .A1(_04226_),
    .S(_03295_),
    .X(_04227_));
 sky130_fd_sc_hd__buf_1 _10068_ (.A(_03292_),
    .X(_04228_));
 sky130_fd_sc_hd__mux2_2 _10069_ (.A0(_04223_),
    .A1(_04227_),
    .S(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_2 _10070_ (.A0(\core.cpuregs[12][0] ),
    .A1(\core.cpuregs[13][0] ),
    .A2(\core.cpuregs[14][0] ),
    .A3(\core.cpuregs[15][0] ),
    .S0(_04218_),
    .S1(_04224_),
    .X(_04230_));
 sky130_fd_sc_hd__mux4_2 _10071_ (.A0(\core.cpuregs[8][0] ),
    .A1(\core.cpuregs[9][0] ),
    .A2(\core.cpuregs[10][0] ),
    .A3(\core.cpuregs[11][0] ),
    .S0(_04218_),
    .S1(_04224_),
    .X(_04231_));
 sky130_fd_sc_hd__mux2_2 _10072_ (.A0(_04230_),
    .A1(_04231_),
    .S(_03295_),
    .X(_04232_));
 sky130_fd_sc_hd__buf_1 _10073_ (.A(_04217_),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_2 _10074_ (.A0(\core.cpuregs[0][0] ),
    .A1(\core.cpuregs[1][0] ),
    .A2(\core.cpuregs[2][0] ),
    .A3(\core.cpuregs[3][0] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04234_));
 sky130_fd_sc_hd__buf_1 _10075_ (.A(_03271_),
    .X(_04235_));
 sky130_fd_sc_hd__buf_1 _10076_ (.A(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__buf_1 _10077_ (.A(_04219_),
    .X(_04237_));
 sky130_fd_sc_hd__mux4_2 _10078_ (.A0(\core.cpuregs[4][0] ),
    .A1(\core.cpuregs[5][0] ),
    .A2(\core.cpuregs[6][0] ),
    .A3(\core.cpuregs[7][0] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__mux2_2 _10079_ (.A0(_04234_),
    .A1(_04238_),
    .S(_03269_),
    .X(_04239_));
 sky130_fd_sc_hd__buf_1 _10080_ (.A(_03309_),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_2 _10081_ (.A0(_04232_),
    .A1(_04239_),
    .S(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__buf_1 _10082_ (.A(_03313_),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_2 _10083_ (.A0(_04229_),
    .A1(_04241_),
    .S(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__buf_1 _10084_ (.A(\core.cpu_state[4] ),
    .X(_04244_));
 sky130_fd_sc_hd__buf_1 _10085_ (.A(_03469_),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_2 _10086_ (.A0(_02475_),
    .A1(_02355_),
    .S(_02099_),
    .X(_04246_));
 sky130_fd_sc_hd__or2_2 _10087_ (.A(_02070_),
    .B(\core.decoded_imm[0] ),
    .X(_04247_));
 sky130_fd_sc_hd__and3_2 _10088_ (.A(_02041_),
    .B(_03415_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__a31o_2 _10089_ (.A1(_04244_),
    .A2(_04245_),
    .A3(_04246_),
    .B1(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__a31o_2 _10090_ (.A1(_03262_),
    .A2(_03265_),
    .A3(_04243_),
    .B1(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__buf_1 _10091_ (.A(_03473_),
    .X(_04251_));
 sky130_fd_sc_hd__mux2_2 _10092_ (.A0(_04250_),
    .A1(_02070_),
    .S(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__buf_1 _10093_ (.A(_04252_),
    .X(_00243_));
 sky130_fd_sc_hd__buf_1 _10094_ (.A(_03339_),
    .X(_04253_));
 sky130_fd_sc_hd__buf_1 _10095_ (.A(_03269_),
    .X(_04254_));
 sky130_fd_sc_hd__buf_1 _10096_ (.A(_03281_),
    .X(_04255_));
 sky130_fd_sc_hd__buf_1 _10097_ (.A(_03278_),
    .X(_04256_));
 sky130_fd_sc_hd__mux4_2 _10098_ (.A0(\core.cpuregs[0][1] ),
    .A1(\core.cpuregs[1][1] ),
    .A2(\core.cpuregs[2][1] ),
    .A3(\core.cpuregs[3][1] ),
    .S0(_04255_),
    .S1(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__or2_2 _10099_ (.A(_04254_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__buf_1 _10100_ (.A(_03289_),
    .X(_04259_));
 sky130_fd_sc_hd__buf_1 _10101_ (.A(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__buf_1 _10102_ (.A(_03271_),
    .X(_04261_));
 sky130_fd_sc_hd__buf_1 _10103_ (.A(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__mux4_2 _10104_ (.A0(\core.cpuregs[4][1] ),
    .A1(\core.cpuregs[5][1] ),
    .A2(\core.cpuregs[6][1] ),
    .A3(\core.cpuregs[7][1] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04263_));
 sky130_fd_sc_hd__or2_2 _10105_ (.A(_04260_),
    .B(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__buf_1 _10106_ (.A(_03266_),
    .X(_04265_));
 sky130_fd_sc_hd__buf_1 _10107_ (.A(_03289_),
    .X(_04266_));
 sky130_fd_sc_hd__buf_1 _10108_ (.A(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__buf_1 _10109_ (.A(_03281_),
    .X(_04268_));
 sky130_fd_sc_hd__mux4_2 _10110_ (.A0(\core.cpuregs[12][1] ),
    .A1(\core.cpuregs[13][1] ),
    .A2(\core.cpuregs[14][1] ),
    .A3(\core.cpuregs[15][1] ),
    .S0(_04268_),
    .S1(_03279_),
    .X(_04269_));
 sky130_fd_sc_hd__mux4_2 _10111_ (.A0(\core.cpuregs[8][1] ),
    .A1(\core.cpuregs[9][1] ),
    .A2(\core.cpuregs[10][1] ),
    .A3(\core.cpuregs[11][1] ),
    .S0(_03281_),
    .S1(_03278_),
    .X(_04270_));
 sky130_fd_sc_hd__or2_2 _10112_ (.A(_03269_),
    .B(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__o211a_2 _10113_ (.A1(_04267_),
    .A2(_04269_),
    .B1(_04271_),
    .C1(_04228_),
    .X(_04272_));
 sky130_fd_sc_hd__a311o_2 _10114_ (.A1(_04240_),
    .A2(_04258_),
    .A3(_04264_),
    .B1(_04265_),
    .C1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__buf_1 _10115_ (.A(_03278_),
    .X(_04274_));
 sky130_fd_sc_hd__mux4_2 _10116_ (.A0(\core.cpuregs[28][1] ),
    .A1(\core.cpuregs[29][1] ),
    .A2(\core.cpuregs[30][1] ),
    .A3(\core.cpuregs[31][1] ),
    .S0(_04268_),
    .S1(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__buf_1 _10117_ (.A(_03283_),
    .X(_04276_));
 sky130_fd_sc_hd__buf_1 _10118_ (.A(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__mux2_2 _10119_ (.A0(\core.cpuregs[24][1] ),
    .A1(\core.cpuregs[25][1] ),
    .S(_03273_),
    .X(_04278_));
 sky130_fd_sc_hd__buf_1 _10120_ (.A(_03271_),
    .X(_04279_));
 sky130_fd_sc_hd__mux2_2 _10121_ (.A0(\core.cpuregs[26][1] ),
    .A1(\core.cpuregs[27][1] ),
    .S(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__buf_1 _10122_ (.A(_03314_),
    .X(_04281_));
 sky130_fd_sc_hd__a21o_2 _10123_ (.A1(_03275_),
    .A2(_04280_),
    .B1(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__a21o_2 _10124_ (.A1(_04277_),
    .A2(_04278_),
    .B1(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__o211a_2 _10125_ (.A1(_04267_),
    .A2(_04275_),
    .B1(_04283_),
    .C1(_04228_),
    .X(_04284_));
 sky130_fd_sc_hd__buf_1 _10126_ (.A(_03275_),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_2 _10127_ (.A0(\core.cpuregs[22][1] ),
    .A1(\core.cpuregs[23][1] ),
    .S(_04268_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_2 _10128_ (.A(_04285_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__mux2_2 _10129_ (.A0(\core.cpuregs[20][1] ),
    .A1(\core.cpuregs[21][1] ),
    .S(_04268_),
    .X(_04288_));
 sky130_fd_sc_hd__a21oi_2 _10130_ (.A1(_04277_),
    .A2(_04288_),
    .B1(_04267_),
    .Y(_04289_));
 sky130_fd_sc_hd__mux4_2 _10131_ (.A0(\core.cpuregs[16][1] ),
    .A1(\core.cpuregs[17][1] ),
    .A2(\core.cpuregs[18][1] ),
    .A3(\core.cpuregs[19][1] ),
    .S0(_04268_),
    .S1(_03279_),
    .X(_04290_));
 sky130_fd_sc_hd__o21ai_2 _10132_ (.A1(_04254_),
    .A2(_04290_),
    .B1(_04240_),
    .Y(_04291_));
 sky130_fd_sc_hd__a21oi_2 _10133_ (.A1(_04287_),
    .A2(_04289_),
    .B1(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__buf_1 _10134_ (.A(_03264_),
    .X(_04293_));
 sky130_fd_sc_hd__o31a_2 _10135_ (.A1(_03313_),
    .A2(_04284_),
    .A3(_04292_),
    .B1(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__a22o_2 _10136_ (.A1(\core.reg_pc[1] ),
    .A2(_04253_),
    .B1(_04273_),
    .B2(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__o21ai_2 _10137_ (.A1(_03414_),
    .A2(_03415_),
    .B1(_02041_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21oi_2 _10138_ (.A1(_03414_),
    .A2(_03415_),
    .B1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__buf_1 _10139_ (.A(_03469_),
    .X(_04298_));
 sky130_fd_sc_hd__mux2_2 _10140_ (.A0(_02070_),
    .A1(_02372_),
    .S(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__a21o_2 _10141_ (.A1(_02388_),
    .A2(_04245_),
    .B1(_02179_),
    .X(_04300_));
 sky130_fd_sc_hd__o211a_2 _10142_ (.A1(_03344_),
    .A2(_04299_),
    .B1(_04300_),
    .C1(_04244_),
    .X(_04301_));
 sky130_fd_sc_hd__a211o_2 _10143_ (.A1(_03262_),
    .A2(_04295_),
    .B1(_04297_),
    .C1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__mux2_2 _10144_ (.A0(_04302_),
    .A1(_02476_),
    .S(_04251_),
    .X(_04303_));
 sky130_fd_sc_hd__buf_1 _10145_ (.A(_04303_),
    .X(_00244_));
 sky130_fd_sc_hd__o21ai_2 _10146_ (.A1(_03418_),
    .A2(_03413_),
    .B1(_03417_),
    .Y(_04304_));
 sky130_fd_sc_hd__o31a_2 _10147_ (.A1(_03418_),
    .A2(_03413_),
    .A3(_03417_),
    .B1(_02042_),
    .X(_04305_));
 sky130_fd_sc_hd__buf_1 _10148_ (.A(_03270_),
    .X(_04306_));
 sky130_fd_sc_hd__buf_1 _10149_ (.A(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__mux4_2 _10150_ (.A0(\core.cpuregs[12][2] ),
    .A1(\core.cpuregs[13][2] ),
    .A2(\core.cpuregs[14][2] ),
    .A3(\core.cpuregs[15][2] ),
    .S0(_04307_),
    .S1(_03274_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_2 _10151_ (.A0(\core.cpuregs[8][2] ),
    .A1(\core.cpuregs[9][2] ),
    .S(_03280_),
    .X(_04309_));
 sky130_fd_sc_hd__mux2_2 _10152_ (.A0(\core.cpuregs[10][2] ),
    .A1(\core.cpuregs[11][2] ),
    .S(_03270_),
    .X(_04310_));
 sky130_fd_sc_hd__a21o_2 _10153_ (.A1(_03277_),
    .A2(_04310_),
    .B1(_03267_),
    .X(_04311_));
 sky130_fd_sc_hd__a21o_2 _10154_ (.A1(_04276_),
    .A2(_04309_),
    .B1(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__o211a_2 _10155_ (.A1(_03294_),
    .A2(_04308_),
    .B1(_04312_),
    .C1(_00008_),
    .X(_04313_));
 sky130_fd_sc_hd__buf_1 _10156_ (.A(_03271_),
    .X(_04314_));
 sky130_fd_sc_hd__buf_1 _10157_ (.A(_00006_),
    .X(_04315_));
 sky130_fd_sc_hd__mux4_2 _10158_ (.A0(\core.cpuregs[0][2] ),
    .A1(\core.cpuregs[1][2] ),
    .A2(\core.cpuregs[2][2] ),
    .A3(\core.cpuregs[3][2] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__buf_1 _10159_ (.A(_03270_),
    .X(_04317_));
 sky130_fd_sc_hd__mux2_2 _10160_ (.A0(\core.cpuregs[4][2] ),
    .A1(\core.cpuregs[5][2] ),
    .S(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_2 _10161_ (.A(_04276_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__mux2_2 _10162_ (.A0(\core.cpuregs[6][2] ),
    .A1(\core.cpuregs[7][2] ),
    .S(_04317_),
    .X(_04320_));
 sky130_fd_sc_hd__nand2_2 _10163_ (.A(_03274_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__a31o_2 _10164_ (.A1(_03314_),
    .A2(_04319_),
    .A3(_04321_),
    .B1(_00008_),
    .X(_04322_));
 sky130_fd_sc_hd__o21ba_2 _10165_ (.A1(_03315_),
    .A2(_04316_),
    .B1_N(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__or3_2 _10166_ (.A(_00009_),
    .B(_04313_),
    .C(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__buf_1 _10167_ (.A(_03314_),
    .X(_04325_));
 sky130_fd_sc_hd__buf_1 _10168_ (.A(_04317_),
    .X(_04326_));
 sky130_fd_sc_hd__mux4_2 _10169_ (.A0(\core.cpuregs[16][2] ),
    .A1(\core.cpuregs[17][2] ),
    .A2(\core.cpuregs[18][2] ),
    .A3(\core.cpuregs[19][2] ),
    .S0(_04326_),
    .S1(_03274_),
    .X(_04327_));
 sky130_fd_sc_hd__buf_1 _10170_ (.A(_03277_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_2 _10171_ (.A0(\core.cpuregs[22][2] ),
    .A1(\core.cpuregs[23][2] ),
    .S(_03280_),
    .X(_04329_));
 sky130_fd_sc_hd__mux2_2 _10172_ (.A0(\core.cpuregs[20][2] ),
    .A1(\core.cpuregs[21][2] ),
    .S(_03270_),
    .X(_04330_));
 sky130_fd_sc_hd__a21o_2 _10173_ (.A1(_03284_),
    .A2(_04330_),
    .B1(_03288_),
    .X(_04331_));
 sky130_fd_sc_hd__a21o_2 _10174_ (.A1(_04328_),
    .A2(_04329_),
    .B1(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__o211a_2 _10175_ (.A1(_04325_),
    .A2(_04327_),
    .B1(_04332_),
    .C1(_03308_),
    .X(_04333_));
 sky130_fd_sc_hd__mux4_2 _10176_ (.A0(\core.cpuregs[24][2] ),
    .A1(\core.cpuregs[25][2] ),
    .A2(\core.cpuregs[26][2] ),
    .A3(\core.cpuregs[27][2] ),
    .S0(_03272_),
    .S1(_03274_),
    .X(_04334_));
 sky130_fd_sc_hd__mux2_2 _10177_ (.A0(\core.cpuregs[30][2] ),
    .A1(\core.cpuregs[31][2] ),
    .S(_03280_),
    .X(_04335_));
 sky130_fd_sc_hd__mux2_2 _10178_ (.A0(\core.cpuregs[28][2] ),
    .A1(\core.cpuregs[29][2] ),
    .S(_03319_),
    .X(_04336_));
 sky130_fd_sc_hd__a21o_2 _10179_ (.A1(_03284_),
    .A2(_04336_),
    .B1(_03288_),
    .X(_04337_));
 sky130_fd_sc_hd__a21o_2 _10180_ (.A1(_04328_),
    .A2(_04335_),
    .B1(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__o211a_2 _10181_ (.A1(_04325_),
    .A2(_04334_),
    .B1(_04338_),
    .C1(_00008_),
    .X(_04339_));
 sky130_fd_sc_hd__or3_2 _10182_ (.A(_03312_),
    .B(_04333_),
    .C(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__a32o_2 _10183_ (.A1(_03264_),
    .A2(_04324_),
    .A3(_04340_),
    .B1(_03339_),
    .B2(_02493_),
    .X(_04341_));
 sky130_fd_sc_hd__and2_2 _10184_ (.A(_03261_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_2 _10185_ (.A0(_02475_),
    .A1(_02375_),
    .S(_04298_),
    .X(_04343_));
 sky130_fd_sc_hd__a21o_2 _10186_ (.A1(_02383_),
    .A2(_04245_),
    .B1(_02179_),
    .X(_04344_));
 sky130_fd_sc_hd__o211a_2 _10187_ (.A1(_03344_),
    .A2(_04343_),
    .B1(_04344_),
    .C1(_04244_),
    .X(_04345_));
 sky130_fd_sc_hd__a211o_2 _10188_ (.A1(_04304_),
    .A2(_04305_),
    .B1(_04342_),
    .C1(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__mux2_2 _10189_ (.A0(_04346_),
    .A1(_02372_),
    .S(_04251_),
    .X(_04347_));
 sky130_fd_sc_hd__buf_1 _10190_ (.A(_04347_),
    .X(_00245_));
 sky130_fd_sc_hd__mux4_2 _10191_ (.A0(\core.cpuregs[8][3] ),
    .A1(\core.cpuregs[9][3] ),
    .A2(\core.cpuregs[10][3] ),
    .A3(\core.cpuregs[11][3] ),
    .S0(_03273_),
    .S1(_03275_),
    .X(_04348_));
 sky130_fd_sc_hd__mux2_2 _10192_ (.A0(\core.cpuregs[14][3] ),
    .A1(\core.cpuregs[15][3] ),
    .S(_03281_),
    .X(_04349_));
 sky130_fd_sc_hd__mux2_2 _10193_ (.A0(\core.cpuregs[12][3] ),
    .A1(\core.cpuregs[13][3] ),
    .S(_03280_),
    .X(_04350_));
 sky130_fd_sc_hd__a21o_2 _10194_ (.A1(_03285_),
    .A2(_04350_),
    .B1(_03289_),
    .X(_04351_));
 sky130_fd_sc_hd__a21o_2 _10195_ (.A1(_03279_),
    .A2(_04349_),
    .B1(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__o211a_2 _10196_ (.A1(_03269_),
    .A2(_04348_),
    .B1(_04352_),
    .C1(_03292_),
    .X(_04353_));
 sky130_fd_sc_hd__mux4_2 _10197_ (.A0(\core.cpuregs[4][3] ),
    .A1(\core.cpuregs[5][3] ),
    .A2(\core.cpuregs[6][3] ),
    .A3(\core.cpuregs[7][3] ),
    .S0(_03297_),
    .S1(_03275_),
    .X(_04354_));
 sky130_fd_sc_hd__mux2_2 _10198_ (.A0(\core.cpuregs[2][3] ),
    .A1(\core.cpuregs[3][3] ),
    .S(_03301_),
    .X(_04355_));
 sky130_fd_sc_hd__mux2_2 _10199_ (.A0(\core.cpuregs[0][3] ),
    .A1(\core.cpuregs[1][3] ),
    .S(_03304_),
    .X(_04356_));
 sky130_fd_sc_hd__a21o_2 _10200_ (.A1(_03285_),
    .A2(_04356_),
    .B1(_03268_),
    .X(_04357_));
 sky130_fd_sc_hd__a21o_2 _10201_ (.A1(_03279_),
    .A2(_04355_),
    .B1(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__o211a_2 _10202_ (.A1(_03295_),
    .A2(_04354_),
    .B1(_04358_),
    .C1(_03309_),
    .X(_04359_));
 sky130_fd_sc_hd__or3_2 _10203_ (.A(_03266_),
    .B(_04353_),
    .C(_04359_),
    .X(_04360_));
 sky130_fd_sc_hd__mux4_2 _10204_ (.A0(\core.cpuregs[16][3] ),
    .A1(\core.cpuregs[17][3] ),
    .A2(\core.cpuregs[18][3] ),
    .A3(\core.cpuregs[19][3] ),
    .S0(_03297_),
    .S1(_03275_),
    .X(_04361_));
 sky130_fd_sc_hd__mux2_2 _10205_ (.A0(\core.cpuregs[22][3] ),
    .A1(\core.cpuregs[23][3] ),
    .S(_03281_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_2 _10206_ (.A0(\core.cpuregs[20][3] ),
    .A1(\core.cpuregs[21][3] ),
    .S(_03320_),
    .X(_04363_));
 sky130_fd_sc_hd__a21o_2 _10207_ (.A1(_03285_),
    .A2(_04363_),
    .B1(_03289_),
    .X(_04364_));
 sky130_fd_sc_hd__a21o_2 _10208_ (.A1(_03279_),
    .A2(_04362_),
    .B1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__o211a_2 _10209_ (.A1(_03316_),
    .A2(_04361_),
    .B1(_04365_),
    .C1(_03309_),
    .X(_04366_));
 sky130_fd_sc_hd__mux4_2 _10210_ (.A0(\core.cpuregs[24][3] ),
    .A1(\core.cpuregs[25][3] ),
    .A2(\core.cpuregs[26][3] ),
    .A3(\core.cpuregs[27][3] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_04367_));
 sky130_fd_sc_hd__mux2_2 _10211_ (.A0(\core.cpuregs[30][3] ),
    .A1(\core.cpuregs[31][3] ),
    .S(_03301_),
    .X(_04368_));
 sky130_fd_sc_hd__mux2_2 _10212_ (.A0(\core.cpuregs[28][3] ),
    .A1(\core.cpuregs[29][3] ),
    .S(_03329_),
    .X(_04369_));
 sky130_fd_sc_hd__a21o_2 _10213_ (.A1(_03285_),
    .A2(_04369_),
    .B1(_03332_),
    .X(_04370_));
 sky130_fd_sc_hd__a21o_2 _10214_ (.A1(_03327_),
    .A2(_04368_),
    .B1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__o211a_2 _10215_ (.A1(_03316_),
    .A2(_04367_),
    .B1(_04371_),
    .C1(_03336_),
    .X(_04372_));
 sky130_fd_sc_hd__or3_2 _10216_ (.A(_03313_),
    .B(_04366_),
    .C(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a32o_2 _10217_ (.A1(_03265_),
    .A2(_04360_),
    .A3(_04373_),
    .B1(_03340_),
    .B2(\core.reg_pc[3] ),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_2 _10218_ (.A0(_02372_),
    .A1(_02355_),
    .S(_04298_),
    .X(_04375_));
 sky130_fd_sc_hd__a21o_2 _10219_ (.A1(_02380_),
    .A2(_04245_),
    .B1(_02179_),
    .X(_04376_));
 sky130_fd_sc_hd__buf_1 _10220_ (.A(\core.cpu_state[4] ),
    .X(_04377_));
 sky130_fd_sc_hd__o211a_2 _10221_ (.A1(_03344_),
    .A2(_04375_),
    .B1(_04376_),
    .C1(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__inv_2 _10222_ (.A(_03412_),
    .Y(_04379_));
 sky130_fd_sc_hd__nand2_2 _10223_ (.A(_03420_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__a21oi_2 _10224_ (.A1(_03419_),
    .A2(_04380_),
    .B1(_02121_),
    .Y(_04381_));
 sky130_fd_sc_hd__o21a_2 _10225_ (.A1(_03419_),
    .A2(_04380_),
    .B1(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__a211o_2 _10226_ (.A1(_03262_),
    .A2(_04374_),
    .B1(_04378_),
    .C1(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__mux2_2 _10227_ (.A0(_04383_),
    .A1(_02375_),
    .S(_04251_),
    .X(_04384_));
 sky130_fd_sc_hd__buf_1 _10228_ (.A(_04384_),
    .X(_00246_));
 sky130_fd_sc_hd__buf_1 _10229_ (.A(_04307_),
    .X(_04385_));
 sky130_fd_sc_hd__mux4_2 _10230_ (.A0(\core.cpuregs[0][4] ),
    .A1(\core.cpuregs[1][4] ),
    .A2(\core.cpuregs[2][4] ),
    .A3(\core.cpuregs[3][4] ),
    .S0(_04385_),
    .S1(_03275_),
    .X(_04386_));
 sky130_fd_sc_hd__buf_1 _10231_ (.A(_03274_),
    .X(_04387_));
 sky130_fd_sc_hd__mux4_2 _10232_ (.A0(\core.cpuregs[4][4] ),
    .A1(\core.cpuregs[5][4] ),
    .A2(\core.cpuregs[6][4] ),
    .A3(\core.cpuregs[7][4] ),
    .S0(_03301_),
    .S1(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__mux4_2 _10233_ (.A0(\core.cpuregs[8][4] ),
    .A1(\core.cpuregs[9][4] ),
    .A2(\core.cpuregs[10][4] ),
    .A3(\core.cpuregs[11][4] ),
    .S0(_03301_),
    .S1(_04387_),
    .X(_04389_));
 sky130_fd_sc_hd__mux4_2 _10234_ (.A0(\core.cpuregs[12][4] ),
    .A1(\core.cpuregs[13][4] ),
    .A2(\core.cpuregs[14][4] ),
    .A3(\core.cpuregs[15][4] ),
    .S0(_03301_),
    .S1(_04387_),
    .X(_04390_));
 sky130_fd_sc_hd__mux4_2 _10235_ (.A0(_04386_),
    .A1(_04388_),
    .A2(_04389_),
    .A3(_04390_),
    .S0(_03269_),
    .S1(_03292_),
    .X(_04391_));
 sky130_fd_sc_hd__or2_2 _10236_ (.A(_04265_),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__mux4_2 _10237_ (.A0(\core.cpuregs[28][4] ),
    .A1(\core.cpuregs[29][4] ),
    .A2(\core.cpuregs[30][4] ),
    .A3(\core.cpuregs[31][4] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_04393_));
 sky130_fd_sc_hd__mux2_2 _10238_ (.A0(\core.cpuregs[24][4] ),
    .A1(\core.cpuregs[25][4] ),
    .S(_03301_),
    .X(_04394_));
 sky130_fd_sc_hd__mux2_2 _10239_ (.A0(\core.cpuregs[26][4] ),
    .A1(\core.cpuregs[27][4] ),
    .S(_03329_),
    .X(_04395_));
 sky130_fd_sc_hd__a21o_2 _10240_ (.A1(_03326_),
    .A2(_04395_),
    .B1(_03268_),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_2 _10241_ (.A1(_04277_),
    .A2(_04394_),
    .B1(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__o211a_2 _10242_ (.A1(_04260_),
    .A2(_04393_),
    .B1(_04397_),
    .C1(_03336_),
    .X(_04398_));
 sky130_fd_sc_hd__buf_1 _10243_ (.A(_04235_),
    .X(_04399_));
 sky130_fd_sc_hd__buf_1 _10244_ (.A(_04219_),
    .X(_04400_));
 sky130_fd_sc_hd__mux4_2 _10245_ (.A0(\core.cpuregs[20][4] ),
    .A1(\core.cpuregs[21][4] ),
    .A2(\core.cpuregs[22][4] ),
    .A3(\core.cpuregs[23][4] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__mux2_2 _10246_ (.A0(\core.cpuregs[18][4] ),
    .A1(\core.cpuregs[19][4] ),
    .S(_03301_),
    .X(_04402_));
 sky130_fd_sc_hd__buf_1 _10247_ (.A(_03283_),
    .X(_04403_));
 sky130_fd_sc_hd__buf_1 _10248_ (.A(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__mux2_2 _10249_ (.A0(\core.cpuregs[16][4] ),
    .A1(\core.cpuregs[17][4] ),
    .S(_04307_),
    .X(_04405_));
 sky130_fd_sc_hd__a21o_2 _10250_ (.A1(_04404_),
    .A2(_04405_),
    .B1(_03268_),
    .X(_04406_));
 sky130_fd_sc_hd__a21o_2 _10251_ (.A1(_03327_),
    .A2(_04402_),
    .B1(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__buf_1 _10252_ (.A(_03308_),
    .X(_04408_));
 sky130_fd_sc_hd__buf_1 _10253_ (.A(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__o211a_2 _10254_ (.A1(_04260_),
    .A2(_04401_),
    .B1(_04407_),
    .C1(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__or3_2 _10255_ (.A(_03313_),
    .B(_04398_),
    .C(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__a32o_2 _10256_ (.A1(_03265_),
    .A2(_04392_),
    .A3(_04411_),
    .B1(_03340_),
    .B2(\core.reg_pc[4] ),
    .X(_04412_));
 sky130_fd_sc_hd__xnor2_2 _10257_ (.A(_03411_),
    .B(_03421_),
    .Y(_04413_));
 sky130_fd_sc_hd__mux4_2 _10258_ (.A0(_02070_),
    .A1(_02375_),
    .A2(_02327_),
    .A3(_02388_),
    .S0(_02178_),
    .S1(_04245_),
    .X(_04414_));
 sky130_fd_sc_hd__a2bb2o_2 _10259_ (.A1_N(_02121_),
    .A2_N(_04413_),
    .B1(_04414_),
    .B2(_02545_),
    .X(_04415_));
 sky130_fd_sc_hd__a31o_2 _10260_ (.A1(_02126_),
    .A2(_02121_),
    .A3(_04412_),
    .B1(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__mux2_2 _10261_ (.A0(_04416_),
    .A1(_02355_),
    .S(_04251_),
    .X(_04417_));
 sky130_fd_sc_hd__buf_1 _10262_ (.A(_04417_),
    .X(_00247_));
 sky130_fd_sc_hd__nor2_2 _10263_ (.A(_03411_),
    .B(_03421_),
    .Y(_04418_));
 sky130_fd_sc_hd__inv_2 _10264_ (.A(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a21oi_2 _10265_ (.A1(_03409_),
    .A2(_04419_),
    .B1(_03408_),
    .Y(_04420_));
 sky130_fd_sc_hd__a31o_2 _10266_ (.A1(_03408_),
    .A2(_03409_),
    .A3(_04419_),
    .B1(_02121_),
    .X(_04421_));
 sky130_fd_sc_hd__mux4_2 _10267_ (.A0(_02475_),
    .A1(_02355_),
    .A2(_02331_),
    .A3(_02383_),
    .S0(_02179_),
    .S1(_04245_),
    .X(_04422_));
 sky130_fd_sc_hd__nand2_2 _10268_ (.A(_02116_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__buf_1 _10269_ (.A(_03262_),
    .X(_04424_));
 sky130_fd_sc_hd__mux4_2 _10270_ (.A0(\core.cpuregs[8][5] ),
    .A1(\core.cpuregs[9][5] ),
    .A2(\core.cpuregs[10][5] ),
    .A3(\core.cpuregs[11][5] ),
    .S0(_03297_),
    .S1(_03275_),
    .X(_04425_));
 sky130_fd_sc_hd__mux2_2 _10271_ (.A0(\core.cpuregs[14][5] ),
    .A1(\core.cpuregs[15][5] ),
    .S(_03281_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_2 _10272_ (.A0(\core.cpuregs[12][5] ),
    .A1(\core.cpuregs[13][5] ),
    .S(_03304_),
    .X(_04427_));
 sky130_fd_sc_hd__a21o_2 _10273_ (.A1(_03285_),
    .A2(_04427_),
    .B1(_03332_),
    .X(_04428_));
 sky130_fd_sc_hd__a21o_2 _10274_ (.A1(_03279_),
    .A2(_04426_),
    .B1(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__o211a_2 _10275_ (.A1(_03316_),
    .A2(_04425_),
    .B1(_04429_),
    .C1(_03336_),
    .X(_04430_));
 sky130_fd_sc_hd__buf_1 _10276_ (.A(_03271_),
    .X(_04431_));
 sky130_fd_sc_hd__buf_1 _10277_ (.A(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__buf_1 _10278_ (.A(_03277_),
    .X(_04433_));
 sky130_fd_sc_hd__buf_1 _10279_ (.A(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__mux4_2 _10280_ (.A0(\core.cpuregs[4][5] ),
    .A1(\core.cpuregs[5][5] ),
    .A2(\core.cpuregs[6][5] ),
    .A3(\core.cpuregs[7][5] ),
    .S0(_04432_),
    .S1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__mux2_2 _10281_ (.A0(\core.cpuregs[2][5] ),
    .A1(\core.cpuregs[3][5] ),
    .S(_03301_),
    .X(_04436_));
 sky130_fd_sc_hd__buf_1 _10282_ (.A(_04306_),
    .X(_04437_));
 sky130_fd_sc_hd__mux2_2 _10283_ (.A0(\core.cpuregs[0][5] ),
    .A1(\core.cpuregs[1][5] ),
    .S(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__a21o_2 _10284_ (.A1(_03285_),
    .A2(_04438_),
    .B1(_03268_),
    .X(_04439_));
 sky130_fd_sc_hd__a21o_2 _10285_ (.A1(_03327_),
    .A2(_04436_),
    .B1(_04439_),
    .X(_04440_));
 sky130_fd_sc_hd__o211a_2 _10286_ (.A1(_04260_),
    .A2(_04435_),
    .B1(_04440_),
    .C1(_04409_),
    .X(_04441_));
 sky130_fd_sc_hd__or3_2 _10287_ (.A(_03266_),
    .B(_04430_),
    .C(_04441_),
    .X(_04442_));
 sky130_fd_sc_hd__mux4_2 _10288_ (.A0(\core.cpuregs[24][5] ),
    .A1(\core.cpuregs[25][5] ),
    .A2(\core.cpuregs[26][5] ),
    .A3(\core.cpuregs[27][5] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_04443_));
 sky130_fd_sc_hd__or2_2 _10289_ (.A(_03316_),
    .B(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__mux2_2 _10290_ (.A0(\core.cpuregs[30][5] ),
    .A1(\core.cpuregs[31][5] ),
    .S(_04268_),
    .X(_04445_));
 sky130_fd_sc_hd__buf_1 _10291_ (.A(_04307_),
    .X(_04446_));
 sky130_fd_sc_hd__mux2_2 _10292_ (.A0(\core.cpuregs[28][5] ),
    .A1(\core.cpuregs[29][5] ),
    .S(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__a21o_2 _10293_ (.A1(_04277_),
    .A2(_04447_),
    .B1(_04266_),
    .X(_04448_));
 sky130_fd_sc_hd__a21o_2 _10294_ (.A1(_04285_),
    .A2(_04445_),
    .B1(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__mux4_2 _10295_ (.A0(\core.cpuregs[20][5] ),
    .A1(\core.cpuregs[21][5] ),
    .A2(\core.cpuregs[22][5] ),
    .A3(\core.cpuregs[23][5] ),
    .S0(_04268_),
    .S1(_03279_),
    .X(_04450_));
 sky130_fd_sc_hd__mux2_2 _10296_ (.A0(\core.cpuregs[16][5] ),
    .A1(\core.cpuregs[17][5] ),
    .S(_03273_),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_2 _10297_ (.A0(\core.cpuregs[18][5] ),
    .A1(\core.cpuregs[19][5] ),
    .S(_03296_),
    .X(_04452_));
 sky130_fd_sc_hd__a21o_2 _10298_ (.A1(_03275_),
    .A2(_04452_),
    .B1(_04325_),
    .X(_04453_));
 sky130_fd_sc_hd__a21o_2 _10299_ (.A1(_04277_),
    .A2(_04451_),
    .B1(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__o211a_2 _10300_ (.A1(_04267_),
    .A2(_04450_),
    .B1(_04454_),
    .C1(_04240_),
    .X(_04455_));
 sky130_fd_sc_hd__a311o_2 _10301_ (.A1(_04228_),
    .A2(_04444_),
    .A3(_04449_),
    .B1(_03313_),
    .C1(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__a32o_2 _10302_ (.A1(_03265_),
    .A2(_04442_),
    .A3(_04456_),
    .B1(_03340_),
    .B2(\core.reg_pc[5] ),
    .X(_04457_));
 sky130_fd_sc_hd__nand2_2 _10303_ (.A(_04424_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__o211ai_2 _10304_ (.A1(_04420_),
    .A2(_04421_),
    .B1(_04423_),
    .C1(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__mux2_2 _10305_ (.A0(_04459_),
    .A1(_02388_),
    .S(_04251_),
    .X(_04460_));
 sky130_fd_sc_hd__buf_1 _10306_ (.A(_04460_),
    .X(_00248_));
 sky130_fd_sc_hd__or2_2 _10307_ (.A(_03408_),
    .B(_04419_),
    .X(_04461_));
 sky130_fd_sc_hd__nand3_2 _10308_ (.A(_03424_),
    .B(_04461_),
    .C(_03431_),
    .Y(_04462_));
 sky130_fd_sc_hd__a21o_2 _10309_ (.A1(_04461_),
    .A2(_03431_),
    .B1(_03424_),
    .X(_04463_));
 sky130_fd_sc_hd__mux4_2 _10310_ (.A0(_02372_),
    .A1(_02388_),
    .A2(_02323_),
    .A3(_02380_),
    .S0(_02178_),
    .S1(_04245_),
    .X(_04464_));
 sky130_fd_sc_hd__a32o_2 _10311_ (.A1(_02041_),
    .A2(_04462_),
    .A3(_04463_),
    .B1(_04464_),
    .B2(_04244_),
    .X(_04465_));
 sky130_fd_sc_hd__mux4_2 _10312_ (.A0(\core.cpuregs[8][6] ),
    .A1(\core.cpuregs[9][6] ),
    .A2(\core.cpuregs[10][6] ),
    .A3(\core.cpuregs[11][6] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04466_));
 sky130_fd_sc_hd__buf_1 _10313_ (.A(_04387_),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_2 _10314_ (.A0(\core.cpuregs[14][6] ),
    .A1(\core.cpuregs[15][6] ),
    .S(_04446_),
    .X(_04468_));
 sky130_fd_sc_hd__buf_1 _10315_ (.A(_04276_),
    .X(_04469_));
 sky130_fd_sc_hd__mux2_2 _10316_ (.A0(\core.cpuregs[12][6] ),
    .A1(\core.cpuregs[13][6] ),
    .S(_03272_),
    .X(_04470_));
 sky130_fd_sc_hd__a21o_2 _10317_ (.A1(_04469_),
    .A2(_04470_),
    .B1(_03294_),
    .X(_04471_));
 sky130_fd_sc_hd__a21o_2 _10318_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__o211a_2 _10319_ (.A1(_04254_),
    .A2(_04466_),
    .B1(_04472_),
    .C1(_04228_),
    .X(_04473_));
 sky130_fd_sc_hd__mux4_2 _10320_ (.A0(\core.cpuregs[4][6] ),
    .A1(\core.cpuregs[5][6] ),
    .A2(\core.cpuregs[6][6] ),
    .A3(\core.cpuregs[7][6] ),
    .S0(_04268_),
    .S1(_04274_),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_2 _10321_ (.A0(\core.cpuregs[2][6] ),
    .A1(\core.cpuregs[3][6] ),
    .S(_03273_),
    .X(_04475_));
 sky130_fd_sc_hd__mux2_2 _10322_ (.A0(\core.cpuregs[0][6] ),
    .A1(\core.cpuregs[1][6] ),
    .S(_04279_),
    .X(_04476_));
 sky130_fd_sc_hd__a21o_2 _10323_ (.A1(_04277_),
    .A2(_04476_),
    .B1(_04281_),
    .X(_04477_));
 sky130_fd_sc_hd__a21o_2 _10324_ (.A1(_04285_),
    .A2(_04475_),
    .B1(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__o211a_2 _10325_ (.A1(_04267_),
    .A2(_04474_),
    .B1(_04478_),
    .C1(_04240_),
    .X(_04479_));
 sky130_fd_sc_hd__or3_2 _10326_ (.A(_04265_),
    .B(_04473_),
    .C(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__mux4_2 _10327_ (.A0(\core.cpuregs[28][6] ),
    .A1(\core.cpuregs[29][6] ),
    .A2(\core.cpuregs[30][6] ),
    .A3(\core.cpuregs[31][6] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04481_));
 sky130_fd_sc_hd__buf_1 _10328_ (.A(_04431_),
    .X(_04482_));
 sky130_fd_sc_hd__mux4_2 _10329_ (.A0(\core.cpuregs[24][6] ),
    .A1(\core.cpuregs[25][6] ),
    .A2(\core.cpuregs[26][6] ),
    .A3(\core.cpuregs[27][6] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04483_));
 sky130_fd_sc_hd__buf_1 _10330_ (.A(_04219_),
    .X(_04484_));
 sky130_fd_sc_hd__mux4_2 _10331_ (.A0(\core.cpuregs[20][6] ),
    .A1(\core.cpuregs[21][6] ),
    .A2(\core.cpuregs[22][6] ),
    .A3(\core.cpuregs[23][6] ),
    .S0(_04399_),
    .S1(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__mux4_2 _10332_ (.A0(\core.cpuregs[16][6] ),
    .A1(\core.cpuregs[17][6] ),
    .A2(\core.cpuregs[18][6] ),
    .A3(\core.cpuregs[19][6] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_04486_));
 sky130_fd_sc_hd__buf_1 _10333_ (.A(_03309_),
    .X(_04487_));
 sky130_fd_sc_hd__mux4_2 _10334_ (.A0(_04481_),
    .A1(_04483_),
    .A2(_04485_),
    .A3(_04486_),
    .S0(_03295_),
    .S1(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__o21a_2 _10335_ (.A1(_04242_),
    .A2(_04488_),
    .B1(_03265_),
    .X(_04489_));
 sky130_fd_sc_hd__nand2_2 _10336_ (.A(_02126_),
    .B(_02121_),
    .Y(_04490_));
 sky130_fd_sc_hd__buf_1 _10337_ (.A(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__a221o_2 _10338_ (.A1(\core.reg_pc[6] ),
    .A2(_03340_),
    .B1(_04480_),
    .B2(_04489_),
    .C1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__o21a_2 _10339_ (.A1(_04424_),
    .A2(_04465_),
    .B1(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__mux2_2 _10340_ (.A0(_04493_),
    .A1(_02383_),
    .S(_04251_),
    .X(_04494_));
 sky130_fd_sc_hd__buf_1 _10341_ (.A(_04494_),
    .X(_00249_));
 sky130_fd_sc_hd__and2_2 _10342_ (.A(_03422_),
    .B(_04463_),
    .X(_04495_));
 sky130_fd_sc_hd__or2_2 _10343_ (.A(_03427_),
    .B(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__nand2_2 _10344_ (.A(_03427_),
    .B(_04495_),
    .Y(_04497_));
 sky130_fd_sc_hd__mux4_2 _10345_ (.A0(_02375_),
    .A1(_02383_),
    .A2(_02336_),
    .A3(_02327_),
    .S0(_02178_),
    .S1(_04245_),
    .X(_04498_));
 sky130_fd_sc_hd__buf_1 _10346_ (.A(_03264_),
    .X(_04499_));
 sky130_fd_sc_hd__buf_1 _10347_ (.A(_00009_),
    .X(_04500_));
 sky130_fd_sc_hd__mux4_2 _10348_ (.A0(\core.cpuregs[8][7] ),
    .A1(\core.cpuregs[9][7] ),
    .A2(\core.cpuregs[10][7] ),
    .A3(\core.cpuregs[11][7] ),
    .S0(_04431_),
    .S1(_03298_),
    .X(_04501_));
 sky130_fd_sc_hd__buf_1 _10349_ (.A(_03277_),
    .X(_04502_));
 sky130_fd_sc_hd__mux2_2 _10350_ (.A0(\core.cpuregs[14][7] ),
    .A1(\core.cpuregs[15][7] ),
    .S(_03320_),
    .X(_04503_));
 sky130_fd_sc_hd__buf_1 _10351_ (.A(_03283_),
    .X(_04504_));
 sky130_fd_sc_hd__mux2_2 _10352_ (.A0(\core.cpuregs[12][7] ),
    .A1(\core.cpuregs[13][7] ),
    .S(_03303_),
    .X(_04505_));
 sky130_fd_sc_hd__a21o_2 _10353_ (.A1(_04504_),
    .A2(_04505_),
    .B1(_03331_),
    .X(_04506_));
 sky130_fd_sc_hd__a21o_2 _10354_ (.A1(_04502_),
    .A2(_04503_),
    .B1(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__buf_1 _10355_ (.A(_00008_),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_2 _10356_ (.A1(_03315_),
    .A2(_04501_),
    .B1(_04507_),
    .C1(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__mux4_2 _10357_ (.A0(\core.cpuregs[4][7] ),
    .A1(\core.cpuregs[5][7] ),
    .A2(\core.cpuregs[6][7] ),
    .A3(\core.cpuregs[7][7] ),
    .S0(_04235_),
    .S1(_04433_),
    .X(_04510_));
 sky130_fd_sc_hd__mux2_2 _10358_ (.A0(\core.cpuregs[2][7] ),
    .A1(\core.cpuregs[3][7] ),
    .S(_03329_),
    .X(_04511_));
 sky130_fd_sc_hd__buf_1 _10359_ (.A(_03283_),
    .X(_04512_));
 sky130_fd_sc_hd__mux2_2 _10360_ (.A0(\core.cpuregs[0][7] ),
    .A1(\core.cpuregs[1][7] ),
    .S(_04306_),
    .X(_04513_));
 sky130_fd_sc_hd__a21o_2 _10361_ (.A1(_04512_),
    .A2(_04513_),
    .B1(_03314_),
    .X(_04514_));
 sky130_fd_sc_hd__a21o_2 _10362_ (.A1(_03326_),
    .A2(_04511_),
    .B1(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__o211a_2 _10363_ (.A1(_04259_),
    .A2(_04510_),
    .B1(_04515_),
    .C1(_04408_),
    .X(_04516_));
 sky130_fd_sc_hd__or3_2 _10364_ (.A(_04500_),
    .B(_04509_),
    .C(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__buf_1 _10365_ (.A(_03312_),
    .X(_04518_));
 sky130_fd_sc_hd__buf_1 _10366_ (.A(_03314_),
    .X(_04519_));
 sky130_fd_sc_hd__mux4_2 _10367_ (.A0(\core.cpuregs[16][7] ),
    .A1(\core.cpuregs[17][7] ),
    .A2(\core.cpuregs[18][7] ),
    .A3(\core.cpuregs[19][7] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04520_));
 sky130_fd_sc_hd__buf_1 _10368_ (.A(_03277_),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_2 _10369_ (.A0(\core.cpuregs[22][7] ),
    .A1(\core.cpuregs[23][7] ),
    .S(_03304_),
    .X(_04522_));
 sky130_fd_sc_hd__buf_1 _10370_ (.A(_03283_),
    .X(_04523_));
 sky130_fd_sc_hd__buf_1 _10371_ (.A(_03270_),
    .X(_04524_));
 sky130_fd_sc_hd__mux2_2 _10372_ (.A0(\core.cpuregs[20][7] ),
    .A1(\core.cpuregs[21][7] ),
    .S(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__buf_1 _10373_ (.A(_03287_),
    .X(_04526_));
 sky130_fd_sc_hd__a21o_2 _10374_ (.A1(_04523_),
    .A2(_04525_),
    .B1(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__a21o_2 _10375_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__buf_1 _10376_ (.A(_03308_),
    .X(_04529_));
 sky130_fd_sc_hd__o211a_2 _10377_ (.A1(_04519_),
    .A2(_04520_),
    .B1(_04528_),
    .C1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__buf_1 _10378_ (.A(_03268_),
    .X(_04531_));
 sky130_fd_sc_hd__mux4_2 _10379_ (.A0(\core.cpuregs[24][7] ),
    .A1(\core.cpuregs[25][7] ),
    .A2(\core.cpuregs[26][7] ),
    .A3(\core.cpuregs[27][7] ),
    .S0(_04261_),
    .S1(_04219_),
    .X(_04532_));
 sky130_fd_sc_hd__buf_1 _10380_ (.A(_03277_),
    .X(_04533_));
 sky130_fd_sc_hd__mux2_2 _10381_ (.A0(\core.cpuregs[30][7] ),
    .A1(\core.cpuregs[31][7] ),
    .S(_04437_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2_2 _10382_ (.A0(\core.cpuregs[28][7] ),
    .A1(\core.cpuregs[29][7] ),
    .S(_04317_),
    .X(_04535_));
 sky130_fd_sc_hd__buf_1 _10383_ (.A(_03287_),
    .X(_04536_));
 sky130_fd_sc_hd__a21o_2 _10384_ (.A1(_04403_),
    .A2(_04535_),
    .B1(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__a21o_2 _10385_ (.A1(_04533_),
    .A2(_04534_),
    .B1(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__o211a_2 _10386_ (.A1(_04531_),
    .A2(_04532_),
    .B1(_04538_),
    .C1(_03292_),
    .X(_04539_));
 sky130_fd_sc_hd__or3_2 _10387_ (.A(_04518_),
    .B(_04530_),
    .C(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__buf_1 _10388_ (.A(_03339_),
    .X(_04541_));
 sky130_fd_sc_hd__a32o_2 _10389_ (.A1(_04499_),
    .A2(_04517_),
    .A3(_04540_),
    .B1(_04541_),
    .B2(\core.reg_pc[7] ),
    .X(_04542_));
 sky130_fd_sc_hd__buf_1 _10390_ (.A(_03261_),
    .X(_04543_));
 sky130_fd_sc_hd__a22o_2 _10391_ (.A1(_04377_),
    .A2(_04498_),
    .B1(_04542_),
    .B2(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__a31o_2 _10392_ (.A1(_02235_),
    .A2(_04496_),
    .A3(_04497_),
    .B1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_2 _10393_ (.A0(_04545_),
    .A1(_02380_),
    .S(_04251_),
    .X(_04546_));
 sky130_fd_sc_hd__buf_1 _10394_ (.A(_04546_),
    .X(_00250_));
 sky130_fd_sc_hd__a21o_2 _10395_ (.A1(_03429_),
    .A2(_03433_),
    .B1(_03436_),
    .X(_04547_));
 sky130_fd_sc_hd__nand3_2 _10396_ (.A(_03436_),
    .B(_03429_),
    .C(_03433_),
    .Y(_04548_));
 sky130_fd_sc_hd__mux4_2 _10397_ (.A0(_02380_),
    .A1(_02355_),
    .A2(_02331_),
    .A3(_02315_),
    .S0(_02099_),
    .S1(_04245_),
    .X(_04549_));
 sky130_fd_sc_hd__a32o_2 _10398_ (.A1(_02041_),
    .A2(_04547_),
    .A3(_04548_),
    .B1(_04549_),
    .B2(_04244_),
    .X(_04550_));
 sky130_fd_sc_hd__mux4_2 _10399_ (.A0(\core.cpuregs[8][8] ),
    .A1(\core.cpuregs[9][8] ),
    .A2(\core.cpuregs[10][8] ),
    .A3(\core.cpuregs[11][8] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04551_));
 sky130_fd_sc_hd__mux2_2 _10400_ (.A0(\core.cpuregs[14][8] ),
    .A1(\core.cpuregs[15][8] ),
    .S(_04446_),
    .X(_04552_));
 sky130_fd_sc_hd__mux2_2 _10401_ (.A0(\core.cpuregs[12][8] ),
    .A1(\core.cpuregs[13][8] ),
    .S(_03272_),
    .X(_04553_));
 sky130_fd_sc_hd__a21o_2 _10402_ (.A1(_04469_),
    .A2(_04553_),
    .B1(_03294_),
    .X(_04554_));
 sky130_fd_sc_hd__a21o_2 _10403_ (.A1(_04467_),
    .A2(_04552_),
    .B1(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__o211a_2 _10404_ (.A1(_04254_),
    .A2(_04551_),
    .B1(_04555_),
    .C1(_04228_),
    .X(_04556_));
 sky130_fd_sc_hd__mux4_2 _10405_ (.A0(\core.cpuregs[4][8] ),
    .A1(\core.cpuregs[5][8] ),
    .A2(\core.cpuregs[6][8] ),
    .A3(\core.cpuregs[7][8] ),
    .S0(_04268_),
    .S1(_04274_),
    .X(_04557_));
 sky130_fd_sc_hd__mux2_2 _10406_ (.A0(\core.cpuregs[2][8] ),
    .A1(\core.cpuregs[3][8] ),
    .S(_03273_),
    .X(_04558_));
 sky130_fd_sc_hd__mux2_2 _10407_ (.A0(\core.cpuregs[0][8] ),
    .A1(\core.cpuregs[1][8] ),
    .S(_04279_),
    .X(_04559_));
 sky130_fd_sc_hd__a21o_2 _10408_ (.A1(_04277_),
    .A2(_04559_),
    .B1(_04281_),
    .X(_04560_));
 sky130_fd_sc_hd__a21o_2 _10409_ (.A1(_04285_),
    .A2(_04558_),
    .B1(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__o211a_2 _10410_ (.A1(_04267_),
    .A2(_04557_),
    .B1(_04561_),
    .C1(_04240_),
    .X(_04562_));
 sky130_fd_sc_hd__or3_2 _10411_ (.A(_04265_),
    .B(_04556_),
    .C(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__mux4_2 _10412_ (.A0(\core.cpuregs[28][8] ),
    .A1(\core.cpuregs[29][8] ),
    .A2(\core.cpuregs[30][8] ),
    .A3(\core.cpuregs[31][8] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04564_));
 sky130_fd_sc_hd__mux4_2 _10413_ (.A0(\core.cpuregs[24][8] ),
    .A1(\core.cpuregs[25][8] ),
    .A2(\core.cpuregs[26][8] ),
    .A3(\core.cpuregs[27][8] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04565_));
 sky130_fd_sc_hd__mux4_2 _10414_ (.A0(\core.cpuregs[20][8] ),
    .A1(\core.cpuregs[21][8] ),
    .A2(\core.cpuregs[22][8] ),
    .A3(\core.cpuregs[23][8] ),
    .S0(_04399_),
    .S1(_04484_),
    .X(_04566_));
 sky130_fd_sc_hd__mux4_2 _10415_ (.A0(\core.cpuregs[16][8] ),
    .A1(\core.cpuregs[17][8] ),
    .A2(\core.cpuregs[18][8] ),
    .A3(\core.cpuregs[19][8] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_04567_));
 sky130_fd_sc_hd__mux4_2 _10416_ (.A0(_04564_),
    .A1(_04565_),
    .A2(_04566_),
    .A3(_04567_),
    .S0(_03295_),
    .S1(_04487_),
    .X(_04568_));
 sky130_fd_sc_hd__o21a_2 _10417_ (.A1(_04242_),
    .A2(_04568_),
    .B1(_03265_),
    .X(_04569_));
 sky130_fd_sc_hd__a221o_2 _10418_ (.A1(\core.reg_pc[8] ),
    .A2(_03340_),
    .B1(_04563_),
    .B2(_04569_),
    .C1(_04491_),
    .X(_04570_));
 sky130_fd_sc_hd__o21a_2 _10419_ (.A1(_04424_),
    .A2(_04550_),
    .B1(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_2 _10420_ (.A0(_04571_),
    .A1(_02327_),
    .S(_04251_),
    .X(_04572_));
 sky130_fd_sc_hd__buf_1 _10421_ (.A(_04572_),
    .X(_00251_));
 sky130_fd_sc_hd__a21o_2 _10422_ (.A1(_03395_),
    .A2(_04547_),
    .B1(_03434_),
    .X(_04573_));
 sky130_fd_sc_hd__nand3_2 _10423_ (.A(_03395_),
    .B(_03434_),
    .C(_04547_),
    .Y(_04574_));
 sky130_fd_sc_hd__buf_1 _10424_ (.A(_02178_),
    .X(_04575_));
 sky130_fd_sc_hd__mux4_2 _10425_ (.A0(_02388_),
    .A1(_02312_),
    .A2(_02327_),
    .A3(_02323_),
    .S0(_04298_),
    .S1(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__mux4_2 _10426_ (.A0(\core.cpuregs[8][9] ),
    .A1(\core.cpuregs[9][9] ),
    .A2(\core.cpuregs[10][9] ),
    .A3(\core.cpuregs[11][9] ),
    .S0(_04431_),
    .S1(_03298_),
    .X(_04577_));
 sky130_fd_sc_hd__mux2_2 _10427_ (.A0(\core.cpuregs[14][9] ),
    .A1(\core.cpuregs[15][9] ),
    .S(_03320_),
    .X(_04578_));
 sky130_fd_sc_hd__mux2_2 _10428_ (.A0(\core.cpuregs[12][9] ),
    .A1(\core.cpuregs[13][9] ),
    .S(_03303_),
    .X(_04579_));
 sky130_fd_sc_hd__a21o_2 _10429_ (.A1(_04504_),
    .A2(_04579_),
    .B1(_03331_),
    .X(_04580_));
 sky130_fd_sc_hd__a21o_2 _10430_ (.A1(_04502_),
    .A2(_04578_),
    .B1(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__o211a_2 _10431_ (.A1(_03315_),
    .A2(_04577_),
    .B1(_04581_),
    .C1(_04508_),
    .X(_04582_));
 sky130_fd_sc_hd__buf_1 _10432_ (.A(_03277_),
    .X(_04583_));
 sky130_fd_sc_hd__mux4_2 _10433_ (.A0(\core.cpuregs[4][9] ),
    .A1(\core.cpuregs[5][9] ),
    .A2(\core.cpuregs[6][9] ),
    .A3(\core.cpuregs[7][9] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__mux2_2 _10434_ (.A0(\core.cpuregs[2][9] ),
    .A1(\core.cpuregs[3][9] ),
    .S(_03329_),
    .X(_04585_));
 sky130_fd_sc_hd__mux2_2 _10435_ (.A0(\core.cpuregs[0][9] ),
    .A1(\core.cpuregs[1][9] ),
    .S(_04306_),
    .X(_04586_));
 sky130_fd_sc_hd__a21o_2 _10436_ (.A1(_04512_),
    .A2(_04586_),
    .B1(_03314_),
    .X(_04587_));
 sky130_fd_sc_hd__a21o_2 _10437_ (.A1(_03326_),
    .A2(_04585_),
    .B1(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__o211a_2 _10438_ (.A1(_04259_),
    .A2(_04584_),
    .B1(_04588_),
    .C1(_04408_),
    .X(_04589_));
 sky130_fd_sc_hd__or3_2 _10439_ (.A(_04500_),
    .B(_04582_),
    .C(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__mux4_2 _10440_ (.A0(\core.cpuregs[16][9] ),
    .A1(\core.cpuregs[17][9] ),
    .A2(\core.cpuregs[18][9] ),
    .A3(\core.cpuregs[19][9] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04591_));
 sky130_fd_sc_hd__buf_1 _10441_ (.A(_03303_),
    .X(_04592_));
 sky130_fd_sc_hd__mux2_2 _10442_ (.A0(\core.cpuregs[22][9] ),
    .A1(\core.cpuregs[23][9] ),
    .S(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__mux2_2 _10443_ (.A0(\core.cpuregs[20][9] ),
    .A1(\core.cpuregs[21][9] ),
    .S(_04524_),
    .X(_04594_));
 sky130_fd_sc_hd__a21o_2 _10444_ (.A1(_04523_),
    .A2(_04594_),
    .B1(_04526_),
    .X(_04595_));
 sky130_fd_sc_hd__a21o_2 _10445_ (.A1(_04521_),
    .A2(_04593_),
    .B1(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__o211a_2 _10446_ (.A1(_04519_),
    .A2(_04591_),
    .B1(_04596_),
    .C1(_04529_),
    .X(_04597_));
 sky130_fd_sc_hd__mux4_2 _10447_ (.A0(\core.cpuregs[24][9] ),
    .A1(\core.cpuregs[25][9] ),
    .A2(\core.cpuregs[26][9] ),
    .A3(\core.cpuregs[27][9] ),
    .S0(_04261_),
    .S1(_04219_),
    .X(_04598_));
 sky130_fd_sc_hd__mux2_2 _10448_ (.A0(\core.cpuregs[30][9] ),
    .A1(\core.cpuregs[31][9] ),
    .S(_04437_),
    .X(_04599_));
 sky130_fd_sc_hd__buf_1 _10449_ (.A(_03270_),
    .X(_04600_));
 sky130_fd_sc_hd__mux2_2 _10450_ (.A0(\core.cpuregs[28][9] ),
    .A1(\core.cpuregs[29][9] ),
    .S(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a21o_2 _10451_ (.A1(_04403_),
    .A2(_04601_),
    .B1(_04536_),
    .X(_04602_));
 sky130_fd_sc_hd__a21o_2 _10452_ (.A1(_04533_),
    .A2(_04599_),
    .B1(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__o211a_2 _10453_ (.A1(_04531_),
    .A2(_04598_),
    .B1(_04603_),
    .C1(_03292_),
    .X(_04604_));
 sky130_fd_sc_hd__or3_2 _10454_ (.A(_04518_),
    .B(_04597_),
    .C(_04604_),
    .X(_04605_));
 sky130_fd_sc_hd__a32o_2 _10455_ (.A1(_04499_),
    .A2(_04590_),
    .A3(_04605_),
    .B1(_04541_),
    .B2(\core.reg_pc[9] ),
    .X(_04606_));
 sky130_fd_sc_hd__a22o_2 _10456_ (.A1(_04377_),
    .A2(_04576_),
    .B1(_04606_),
    .B2(_04543_),
    .X(_04607_));
 sky130_fd_sc_hd__a31o_2 _10457_ (.A1(_02235_),
    .A2(_04573_),
    .A3(_04574_),
    .B1(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__mux2_2 _10458_ (.A0(_04608_),
    .A1(_02331_),
    .S(_04251_),
    .X(_04609_));
 sky130_fd_sc_hd__buf_1 _10459_ (.A(_04609_),
    .X(_00252_));
 sky130_fd_sc_hd__nand2_2 _10460_ (.A(_03391_),
    .B(_03392_),
    .Y(_04610_));
 sky130_fd_sc_hd__o21a_2 _10461_ (.A1(_03434_),
    .A2(_04547_),
    .B1(_03397_),
    .X(_04611_));
 sky130_fd_sc_hd__xor2_2 _10462_ (.A(_04610_),
    .B(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__buf_1 _10463_ (.A(_03342_),
    .X(_04613_));
 sky130_fd_sc_hd__mux2_2 _10464_ (.A0(_02336_),
    .A1(_02331_),
    .S(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__mux2_2 _10465_ (.A0(_02383_),
    .A1(_02306_),
    .S(_03469_),
    .X(_04615_));
 sky130_fd_sc_hd__mux2_2 _10466_ (.A0(_04614_),
    .A1(_04615_),
    .S(_03344_),
    .X(_04616_));
 sky130_fd_sc_hd__a22o_2 _10467_ (.A1(_02042_),
    .A2(_04612_),
    .B1(_04616_),
    .B2(_04244_),
    .X(_04617_));
 sky130_fd_sc_hd__mux4_2 _10468_ (.A0(\core.cpuregs[8][10] ),
    .A1(\core.cpuregs[9][10] ),
    .A2(\core.cpuregs[10][10] ),
    .A3(\core.cpuregs[11][10] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04618_));
 sky130_fd_sc_hd__mux2_2 _10469_ (.A0(\core.cpuregs[14][10] ),
    .A1(\core.cpuregs[15][10] ),
    .S(_04446_),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_2 _10470_ (.A0(\core.cpuregs[12][10] ),
    .A1(\core.cpuregs[13][10] ),
    .S(_03272_),
    .X(_04620_));
 sky130_fd_sc_hd__a21o_2 _10471_ (.A1(_04469_),
    .A2(_04620_),
    .B1(_03294_),
    .X(_04621_));
 sky130_fd_sc_hd__a21o_2 _10472_ (.A1(_04467_),
    .A2(_04619_),
    .B1(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__o211a_2 _10473_ (.A1(_04254_),
    .A2(_04618_),
    .B1(_04622_),
    .C1(_04228_),
    .X(_04623_));
 sky130_fd_sc_hd__mux4_2 _10474_ (.A0(\core.cpuregs[4][10] ),
    .A1(\core.cpuregs[5][10] ),
    .A2(\core.cpuregs[6][10] ),
    .A3(\core.cpuregs[7][10] ),
    .S0(_04268_),
    .S1(_04274_),
    .X(_04624_));
 sky130_fd_sc_hd__mux2_2 _10475_ (.A0(\core.cpuregs[2][10] ),
    .A1(\core.cpuregs[3][10] ),
    .S(_03273_),
    .X(_04625_));
 sky130_fd_sc_hd__mux2_2 _10476_ (.A0(\core.cpuregs[0][10] ),
    .A1(\core.cpuregs[1][10] ),
    .S(_04279_),
    .X(_04626_));
 sky130_fd_sc_hd__a21o_2 _10477_ (.A1(_04277_),
    .A2(_04626_),
    .B1(_04281_),
    .X(_04627_));
 sky130_fd_sc_hd__a21o_2 _10478_ (.A1(_04285_),
    .A2(_04625_),
    .B1(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__o211a_2 _10479_ (.A1(_04267_),
    .A2(_04624_),
    .B1(_04628_),
    .C1(_04240_),
    .X(_04629_));
 sky130_fd_sc_hd__or3_2 _10480_ (.A(_04265_),
    .B(_04623_),
    .C(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__mux4_2 _10481_ (.A0(\core.cpuregs[28][10] ),
    .A1(\core.cpuregs[29][10] ),
    .A2(\core.cpuregs[30][10] ),
    .A3(\core.cpuregs[31][10] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04631_));
 sky130_fd_sc_hd__mux4_2 _10482_ (.A0(\core.cpuregs[24][10] ),
    .A1(\core.cpuregs[25][10] ),
    .A2(\core.cpuregs[26][10] ),
    .A3(\core.cpuregs[27][10] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04632_));
 sky130_fd_sc_hd__mux4_2 _10483_ (.A0(\core.cpuregs[20][10] ),
    .A1(\core.cpuregs[21][10] ),
    .A2(\core.cpuregs[22][10] ),
    .A3(\core.cpuregs[23][10] ),
    .S0(_04399_),
    .S1(_04484_),
    .X(_04633_));
 sky130_fd_sc_hd__mux4_2 _10484_ (.A0(\core.cpuregs[16][10] ),
    .A1(\core.cpuregs[17][10] ),
    .A2(\core.cpuregs[18][10] ),
    .A3(\core.cpuregs[19][10] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_04634_));
 sky130_fd_sc_hd__mux4_2 _10485_ (.A0(_04631_),
    .A1(_04632_),
    .A2(_04633_),
    .A3(_04634_),
    .S0(_03295_),
    .S1(_04487_),
    .X(_04635_));
 sky130_fd_sc_hd__o21a_2 _10486_ (.A1(_04242_),
    .A2(_04635_),
    .B1(_03265_),
    .X(_04636_));
 sky130_fd_sc_hd__a221o_2 _10487_ (.A1(\core.reg_pc[10] ),
    .A2(_03340_),
    .B1(_04630_),
    .B2(_04636_),
    .C1(_04491_),
    .X(_04637_));
 sky130_fd_sc_hd__o21a_2 _10488_ (.A1(_04424_),
    .A2(_04617_),
    .B1(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__buf_1 _10489_ (.A(_03473_),
    .X(_04639_));
 sky130_fd_sc_hd__mux2_2 _10490_ (.A0(_04638_),
    .A1(_02323_),
    .S(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__buf_1 _10491_ (.A(_04640_),
    .X(_00253_));
 sky130_fd_sc_hd__o21ai_2 _10492_ (.A1(_04610_),
    .A2(_04611_),
    .B1(_03391_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_2 _10493_ (.A(_03390_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__or2_2 _10494_ (.A(_03390_),
    .B(_04641_),
    .X(_04643_));
 sky130_fd_sc_hd__mux4_2 _10495_ (.A0(_02380_),
    .A1(_02345_),
    .A2(_02323_),
    .A3(_02315_),
    .S0(_04298_),
    .S1(_04575_),
    .X(_04644_));
 sky130_fd_sc_hd__mux4_2 _10496_ (.A0(\core.cpuregs[8][11] ),
    .A1(\core.cpuregs[9][11] ),
    .A2(\core.cpuregs[10][11] ),
    .A3(\core.cpuregs[11][11] ),
    .S0(_04431_),
    .S1(_03298_),
    .X(_04645_));
 sky130_fd_sc_hd__mux2_2 _10497_ (.A0(\core.cpuregs[14][11] ),
    .A1(\core.cpuregs[15][11] ),
    .S(_03320_),
    .X(_04646_));
 sky130_fd_sc_hd__mux2_2 _10498_ (.A0(\core.cpuregs[12][11] ),
    .A1(\core.cpuregs[13][11] ),
    .S(_03303_),
    .X(_04647_));
 sky130_fd_sc_hd__a21o_2 _10499_ (.A1(_04504_),
    .A2(_04647_),
    .B1(_03331_),
    .X(_04648_));
 sky130_fd_sc_hd__a21o_2 _10500_ (.A1(_04502_),
    .A2(_04646_),
    .B1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__o211a_2 _10501_ (.A1(_03315_),
    .A2(_04645_),
    .B1(_04649_),
    .C1(_04508_),
    .X(_04650_));
 sky130_fd_sc_hd__mux4_2 _10502_ (.A0(\core.cpuregs[4][11] ),
    .A1(\core.cpuregs[5][11] ),
    .A2(\core.cpuregs[6][11] ),
    .A3(\core.cpuregs[7][11] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_04651_));
 sky130_fd_sc_hd__mux2_2 _10503_ (.A0(\core.cpuregs[2][11] ),
    .A1(\core.cpuregs[3][11] ),
    .S(_03329_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_2 _10504_ (.A0(\core.cpuregs[0][11] ),
    .A1(\core.cpuregs[1][11] ),
    .S(_04306_),
    .X(_04653_));
 sky130_fd_sc_hd__a21o_2 _10505_ (.A1(_04512_),
    .A2(_04653_),
    .B1(_03314_),
    .X(_04654_));
 sky130_fd_sc_hd__a21o_2 _10506_ (.A1(_03326_),
    .A2(_04652_),
    .B1(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__o211a_2 _10507_ (.A1(_04259_),
    .A2(_04651_),
    .B1(_04655_),
    .C1(_04408_),
    .X(_04656_));
 sky130_fd_sc_hd__or3_2 _10508_ (.A(_04500_),
    .B(_04650_),
    .C(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__mux4_2 _10509_ (.A0(\core.cpuregs[16][11] ),
    .A1(\core.cpuregs[17][11] ),
    .A2(\core.cpuregs[18][11] ),
    .A3(\core.cpuregs[19][11] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_2 _10510_ (.A0(\core.cpuregs[22][11] ),
    .A1(\core.cpuregs[23][11] ),
    .S(_04592_),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_2 _10511_ (.A0(\core.cpuregs[20][11] ),
    .A1(\core.cpuregs[21][11] ),
    .S(_04524_),
    .X(_04660_));
 sky130_fd_sc_hd__a21o_2 _10512_ (.A1(_04523_),
    .A2(_04660_),
    .B1(_04526_),
    .X(_04661_));
 sky130_fd_sc_hd__a21o_2 _10513_ (.A1(_04521_),
    .A2(_04659_),
    .B1(_04661_),
    .X(_04662_));
 sky130_fd_sc_hd__o211a_2 _10514_ (.A1(_04519_),
    .A2(_04658_),
    .B1(_04662_),
    .C1(_04529_),
    .X(_04663_));
 sky130_fd_sc_hd__mux4_2 _10515_ (.A0(\core.cpuregs[24][11] ),
    .A1(\core.cpuregs[25][11] ),
    .A2(\core.cpuregs[26][11] ),
    .A3(\core.cpuregs[27][11] ),
    .S0(_04261_),
    .S1(_04219_),
    .X(_04664_));
 sky130_fd_sc_hd__mux2_2 _10516_ (.A0(\core.cpuregs[30][11] ),
    .A1(\core.cpuregs[31][11] ),
    .S(_04437_),
    .X(_04665_));
 sky130_fd_sc_hd__mux2_2 _10517_ (.A0(\core.cpuregs[28][11] ),
    .A1(\core.cpuregs[29][11] ),
    .S(_04600_),
    .X(_04666_));
 sky130_fd_sc_hd__a21o_2 _10518_ (.A1(_04403_),
    .A2(_04666_),
    .B1(_04536_),
    .X(_04667_));
 sky130_fd_sc_hd__a21o_2 _10519_ (.A1(_04533_),
    .A2(_04665_),
    .B1(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__o211a_2 _10520_ (.A1(_04531_),
    .A2(_04664_),
    .B1(_04668_),
    .C1(_03335_),
    .X(_04669_));
 sky130_fd_sc_hd__or3_2 _10521_ (.A(_04518_),
    .B(_04663_),
    .C(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__a32o_2 _10522_ (.A1(_04499_),
    .A2(_04657_),
    .A3(_04670_),
    .B1(_04541_),
    .B2(\core.reg_pc[11] ),
    .X(_04671_));
 sky130_fd_sc_hd__a22o_2 _10523_ (.A1(_04377_),
    .A2(_04644_),
    .B1(_04671_),
    .B2(_04543_),
    .X(_04672_));
 sky130_fd_sc_hd__a31o_2 _10524_ (.A1(_02235_),
    .A2(_04642_),
    .A3(_04643_),
    .B1(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_2 _10525_ (.A0(_04673_),
    .A1(_02336_),
    .S(_04639_),
    .X(_04674_));
 sky130_fd_sc_hd__buf_1 _10526_ (.A(_04674_),
    .X(_00254_));
 sky130_fd_sc_hd__or3_2 _10527_ (.A(_03393_),
    .B(_03434_),
    .C(_04547_),
    .X(_04675_));
 sky130_fd_sc_hd__a21o_2 _10528_ (.A1(_03400_),
    .A2(_04675_),
    .B1(_03388_),
    .X(_04676_));
 sky130_fd_sc_hd__a31oi_2 _10529_ (.A1(_03388_),
    .A2(_03400_),
    .A3(_04675_),
    .B1(_02121_),
    .Y(_04677_));
 sky130_fd_sc_hd__mux2_2 _10530_ (.A0(_02312_),
    .A1(_02336_),
    .S(_04613_),
    .X(_04678_));
 sky130_fd_sc_hd__mux2_2 _10531_ (.A0(_02327_),
    .A1(_02291_),
    .S(_03469_),
    .X(_04679_));
 sky130_fd_sc_hd__mux2_2 _10532_ (.A0(_04678_),
    .A1(_04679_),
    .S(_03344_),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_2 _10533_ (.A1(_04676_),
    .A2(_04677_),
    .B1(_04680_),
    .B2(_04377_),
    .X(_04681_));
 sky130_fd_sc_hd__mux4_2 _10534_ (.A0(\core.cpuregs[8][12] ),
    .A1(\core.cpuregs[9][12] ),
    .A2(\core.cpuregs[10][12] ),
    .A3(\core.cpuregs[11][12] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04682_));
 sky130_fd_sc_hd__mux2_2 _10535_ (.A0(\core.cpuregs[14][12] ),
    .A1(\core.cpuregs[15][12] ),
    .S(_04385_),
    .X(_04683_));
 sky130_fd_sc_hd__mux2_2 _10536_ (.A0(\core.cpuregs[12][12] ),
    .A1(\core.cpuregs[13][12] ),
    .S(_03272_),
    .X(_04684_));
 sky130_fd_sc_hd__a21o_2 _10537_ (.A1(_04404_),
    .A2(_04684_),
    .B1(_03294_),
    .X(_04685_));
 sky130_fd_sc_hd__a21o_2 _10538_ (.A1(_04467_),
    .A2(_04683_),
    .B1(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__o211a_2 _10539_ (.A1(_04254_),
    .A2(_04682_),
    .B1(_04686_),
    .C1(_04228_),
    .X(_04687_));
 sky130_fd_sc_hd__mux4_2 _10540_ (.A0(\core.cpuregs[4][12] ),
    .A1(\core.cpuregs[5][12] ),
    .A2(\core.cpuregs[6][12] ),
    .A3(\core.cpuregs[7][12] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_04688_));
 sky130_fd_sc_hd__mux2_2 _10541_ (.A0(\core.cpuregs[2][12] ),
    .A1(\core.cpuregs[3][12] ),
    .S(_03273_),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_2 _10542_ (.A0(\core.cpuregs[0][12] ),
    .A1(\core.cpuregs[1][12] ),
    .S(_04279_),
    .X(_04690_));
 sky130_fd_sc_hd__a21o_2 _10543_ (.A1(_04277_),
    .A2(_04690_),
    .B1(_04281_),
    .X(_04691_));
 sky130_fd_sc_hd__a21o_2 _10544_ (.A1(_04285_),
    .A2(_04689_),
    .B1(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__o211a_2 _10545_ (.A1(_04267_),
    .A2(_04688_),
    .B1(_04692_),
    .C1(_04240_),
    .X(_04693_));
 sky130_fd_sc_hd__or3_2 _10546_ (.A(_04265_),
    .B(_04687_),
    .C(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__mux4_2 _10547_ (.A0(\core.cpuregs[28][12] ),
    .A1(\core.cpuregs[29][12] ),
    .A2(\core.cpuregs[30][12] ),
    .A3(\core.cpuregs[31][12] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04695_));
 sky130_fd_sc_hd__mux4_2 _10548_ (.A0(\core.cpuregs[24][12] ),
    .A1(\core.cpuregs[25][12] ),
    .A2(\core.cpuregs[26][12] ),
    .A3(\core.cpuregs[27][12] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04696_));
 sky130_fd_sc_hd__mux4_2 _10549_ (.A0(\core.cpuregs[20][12] ),
    .A1(\core.cpuregs[21][12] ),
    .A2(\core.cpuregs[22][12] ),
    .A3(\core.cpuregs[23][12] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_04697_));
 sky130_fd_sc_hd__mux4_2 _10550_ (.A0(\core.cpuregs[16][12] ),
    .A1(\core.cpuregs[17][12] ),
    .A2(\core.cpuregs[18][12] ),
    .A3(\core.cpuregs[19][12] ),
    .S0(_04236_),
    .S1(_04400_),
    .X(_04698_));
 sky130_fd_sc_hd__mux4_2 _10551_ (.A0(_04695_),
    .A1(_04696_),
    .A2(_04697_),
    .A3(_04698_),
    .S0(_03295_),
    .S1(_04487_),
    .X(_04699_));
 sky130_fd_sc_hd__o21a_2 _10552_ (.A1(_04242_),
    .A2(_04699_),
    .B1(_03265_),
    .X(_04700_));
 sky130_fd_sc_hd__a221o_2 _10553_ (.A1(\core.reg_pc[12] ),
    .A2(_03340_),
    .B1(_04694_),
    .B2(_04700_),
    .C1(_04491_),
    .X(_04701_));
 sky130_fd_sc_hd__o21a_2 _10554_ (.A1(_04424_),
    .A2(_04681_),
    .B1(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__mux2_2 _10555_ (.A0(_04702_),
    .A1(_02315_),
    .S(_04639_),
    .X(_04703_));
 sky130_fd_sc_hd__buf_1 _10556_ (.A(_04703_),
    .X(_00255_));
 sky130_fd_sc_hd__a21o_2 _10557_ (.A1(_03386_),
    .A2(_04676_),
    .B1(_03385_),
    .X(_04704_));
 sky130_fd_sc_hd__nand3_2 _10558_ (.A(_03385_),
    .B(_03386_),
    .C(_04676_),
    .Y(_04705_));
 sky130_fd_sc_hd__mux4_2 _10559_ (.A0(_02306_),
    .A1(_02315_),
    .A2(_02293_),
    .A3(_02331_),
    .S0(_03343_),
    .S1(_02099_),
    .X(_04706_));
 sky130_fd_sc_hd__mux4_2 _10560_ (.A0(\core.cpuregs[8][13] ),
    .A1(\core.cpuregs[9][13] ),
    .A2(\core.cpuregs[10][13] ),
    .A3(\core.cpuregs[11][13] ),
    .S0(_03296_),
    .S1(_03298_),
    .X(_04707_));
 sky130_fd_sc_hd__mux2_2 _10561_ (.A0(\core.cpuregs[14][13] ),
    .A1(\core.cpuregs[15][13] ),
    .S(_03320_),
    .X(_04708_));
 sky130_fd_sc_hd__mux2_2 _10562_ (.A0(\core.cpuregs[12][13] ),
    .A1(\core.cpuregs[13][13] ),
    .S(_03319_),
    .X(_04709_));
 sky130_fd_sc_hd__a21o_2 _10563_ (.A1(_04504_),
    .A2(_04709_),
    .B1(_03331_),
    .X(_04710_));
 sky130_fd_sc_hd__a21o_2 _10564_ (.A1(_04328_),
    .A2(_04708_),
    .B1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__o211a_2 _10565_ (.A1(_03315_),
    .A2(_04707_),
    .B1(_04711_),
    .C1(_04508_),
    .X(_04712_));
 sky130_fd_sc_hd__mux4_2 _10566_ (.A0(\core.cpuregs[4][13] ),
    .A1(\core.cpuregs[5][13] ),
    .A2(\core.cpuregs[6][13] ),
    .A3(\core.cpuregs[7][13] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_04713_));
 sky130_fd_sc_hd__mux2_2 _10567_ (.A0(\core.cpuregs[2][13] ),
    .A1(\core.cpuregs[3][13] ),
    .S(_03329_),
    .X(_04714_));
 sky130_fd_sc_hd__mux2_2 _10568_ (.A0(\core.cpuregs[0][13] ),
    .A1(\core.cpuregs[1][13] ),
    .S(_04306_),
    .X(_04715_));
 sky130_fd_sc_hd__a21o_2 _10569_ (.A1(_04512_),
    .A2(_04715_),
    .B1(_03267_),
    .X(_04716_));
 sky130_fd_sc_hd__a21o_2 _10570_ (.A1(_03326_),
    .A2(_04714_),
    .B1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__o211a_2 _10571_ (.A1(_04259_),
    .A2(_04713_),
    .B1(_04717_),
    .C1(_04408_),
    .X(_04718_));
 sky130_fd_sc_hd__or3_2 _10572_ (.A(_04500_),
    .B(_04712_),
    .C(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__mux4_2 _10573_ (.A0(\core.cpuregs[16][13] ),
    .A1(\core.cpuregs[17][13] ),
    .A2(\core.cpuregs[18][13] ),
    .A3(\core.cpuregs[19][13] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_2 _10574_ (.A0(\core.cpuregs[22][13] ),
    .A1(\core.cpuregs[23][13] ),
    .S(_04592_),
    .X(_04721_));
 sky130_fd_sc_hd__mux2_2 _10575_ (.A0(\core.cpuregs[20][13] ),
    .A1(\core.cpuregs[21][13] ),
    .S(_04524_),
    .X(_04722_));
 sky130_fd_sc_hd__a21o_2 _10576_ (.A1(_04523_),
    .A2(_04722_),
    .B1(_04526_),
    .X(_04723_));
 sky130_fd_sc_hd__a21o_2 _10577_ (.A1(_04521_),
    .A2(_04721_),
    .B1(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__o211a_2 _10578_ (.A1(_04519_),
    .A2(_04720_),
    .B1(_04724_),
    .C1(_04529_),
    .X(_04725_));
 sky130_fd_sc_hd__mux4_2 _10579_ (.A0(\core.cpuregs[24][13] ),
    .A1(\core.cpuregs[25][13] ),
    .A2(\core.cpuregs[26][13] ),
    .A3(\core.cpuregs[27][13] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_2 _10580_ (.A0(\core.cpuregs[30][13] ),
    .A1(\core.cpuregs[31][13] ),
    .S(_04437_),
    .X(_04727_));
 sky130_fd_sc_hd__mux2_2 _10581_ (.A0(\core.cpuregs[28][13] ),
    .A1(\core.cpuregs[29][13] ),
    .S(_04600_),
    .X(_04728_));
 sky130_fd_sc_hd__a21o_2 _10582_ (.A1(_04403_),
    .A2(_04728_),
    .B1(_04536_),
    .X(_04729_));
 sky130_fd_sc_hd__a21o_2 _10583_ (.A1(_04533_),
    .A2(_04727_),
    .B1(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__o211a_2 _10584_ (.A1(_04531_),
    .A2(_04726_),
    .B1(_04730_),
    .C1(_03335_),
    .X(_04731_));
 sky130_fd_sc_hd__or3_2 _10585_ (.A(_04518_),
    .B(_04725_),
    .C(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__a32o_2 _10586_ (.A1(_04499_),
    .A2(_04719_),
    .A3(_04732_),
    .B1(_04541_),
    .B2(\core.reg_pc[13] ),
    .X(_04733_));
 sky130_fd_sc_hd__a22o_2 _10587_ (.A1(_02545_),
    .A2(_04706_),
    .B1(_04733_),
    .B2(_04543_),
    .X(_04734_));
 sky130_fd_sc_hd__a31o_2 _10588_ (.A1(_02235_),
    .A2(_04704_),
    .A3(_04705_),
    .B1(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_2 _10589_ (.A0(_04735_),
    .A1(_02312_),
    .S(_04639_),
    .X(_04736_));
 sky130_fd_sc_hd__buf_1 _10590_ (.A(_04736_),
    .X(_00256_));
 sky130_fd_sc_hd__a31o_2 _10591_ (.A1(_03384_),
    .A2(_03386_),
    .A3(_04676_),
    .B1(_03383_),
    .X(_04737_));
 sky130_fd_sc_hd__nand2_2 _10592_ (.A(_03439_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__o21a_2 _10593_ (.A1(_03439_),
    .A2(_04737_),
    .B1(_02041_),
    .X(_04739_));
 sky130_fd_sc_hd__mux4_2 _10594_ (.A0(_02345_),
    .A1(_02312_),
    .A2(_02298_),
    .A3(_02323_),
    .S0(_03343_),
    .S1(_03344_),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_2 _10595_ (.A1(_04738_),
    .A2(_04739_),
    .B1(_04740_),
    .B2(_04377_),
    .X(_04741_));
 sky130_fd_sc_hd__mux4_2 _10596_ (.A0(\core.cpuregs[8][14] ),
    .A1(\core.cpuregs[9][14] ),
    .A2(\core.cpuregs[10][14] ),
    .A3(\core.cpuregs[11][14] ),
    .S0(_04262_),
    .S1(_04256_),
    .X(_04742_));
 sky130_fd_sc_hd__mux2_2 _10597_ (.A0(\core.cpuregs[14][14] ),
    .A1(\core.cpuregs[15][14] ),
    .S(_04385_),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_2 _10598_ (.A0(\core.cpuregs[12][14] ),
    .A1(\core.cpuregs[13][14] ),
    .S(_03272_),
    .X(_04744_));
 sky130_fd_sc_hd__a21o_2 _10599_ (.A1(_04404_),
    .A2(_04744_),
    .B1(_03294_),
    .X(_04745_));
 sky130_fd_sc_hd__a21o_2 _10600_ (.A1(_04467_),
    .A2(_04743_),
    .B1(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__o211a_2 _10601_ (.A1(_04254_),
    .A2(_04742_),
    .B1(_04746_),
    .C1(_04228_),
    .X(_04747_));
 sky130_fd_sc_hd__mux4_2 _10602_ (.A0(\core.cpuregs[4][14] ),
    .A1(\core.cpuregs[5][14] ),
    .A2(\core.cpuregs[6][14] ),
    .A3(\core.cpuregs[7][14] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_04748_));
 sky130_fd_sc_hd__mux2_2 _10603_ (.A0(\core.cpuregs[2][14] ),
    .A1(\core.cpuregs[3][14] ),
    .S(_03273_),
    .X(_04749_));
 sky130_fd_sc_hd__mux2_2 _10604_ (.A0(\core.cpuregs[0][14] ),
    .A1(\core.cpuregs[1][14] ),
    .S(_04279_),
    .X(_04750_));
 sky130_fd_sc_hd__a21o_2 _10605_ (.A1(_04277_),
    .A2(_04750_),
    .B1(_04281_),
    .X(_04751_));
 sky130_fd_sc_hd__a21o_2 _10606_ (.A1(_04285_),
    .A2(_04749_),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__o211a_2 _10607_ (.A1(_04267_),
    .A2(_04748_),
    .B1(_04752_),
    .C1(_04240_),
    .X(_04753_));
 sky130_fd_sc_hd__or3_2 _10608_ (.A(_04265_),
    .B(_04747_),
    .C(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__mux4_2 _10609_ (.A0(\core.cpuregs[28][14] ),
    .A1(\core.cpuregs[29][14] ),
    .A2(\core.cpuregs[30][14] ),
    .A3(\core.cpuregs[31][14] ),
    .S0(_04233_),
    .S1(_04224_),
    .X(_04755_));
 sky130_fd_sc_hd__mux4_2 _10610_ (.A0(\core.cpuregs[24][14] ),
    .A1(\core.cpuregs[25][14] ),
    .A2(\core.cpuregs[26][14] ),
    .A3(\core.cpuregs[27][14] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04756_));
 sky130_fd_sc_hd__mux4_2 _10611_ (.A0(\core.cpuregs[20][14] ),
    .A1(\core.cpuregs[21][14] ),
    .A2(\core.cpuregs[22][14] ),
    .A3(\core.cpuregs[23][14] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_04757_));
 sky130_fd_sc_hd__mux4_2 _10612_ (.A0(\core.cpuregs[16][14] ),
    .A1(\core.cpuregs[17][14] ),
    .A2(\core.cpuregs[18][14] ),
    .A3(\core.cpuregs[19][14] ),
    .S0(_04236_),
    .S1(_04400_),
    .X(_04758_));
 sky130_fd_sc_hd__mux4_2 _10613_ (.A0(_04755_),
    .A1(_04756_),
    .A2(_04757_),
    .A3(_04758_),
    .S0(_03295_),
    .S1(_04409_),
    .X(_04759_));
 sky130_fd_sc_hd__o21a_2 _10614_ (.A1(_04242_),
    .A2(_04759_),
    .B1(_03265_),
    .X(_04760_));
 sky130_fd_sc_hd__a221o_2 _10615_ (.A1(\core.reg_pc[14] ),
    .A2(_03340_),
    .B1(_04754_),
    .B2(_04760_),
    .C1(_04491_),
    .X(_04761_));
 sky130_fd_sc_hd__o21a_2 _10616_ (.A1(_04424_),
    .A2(_04741_),
    .B1(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__mux2_2 _10617_ (.A0(_04762_),
    .A1(_02306_),
    .S(_04639_),
    .X(_04763_));
 sky130_fd_sc_hd__buf_1 _10618_ (.A(_04763_),
    .X(_00257_));
 sky130_fd_sc_hd__o21ai_2 _10619_ (.A1(_03439_),
    .A2(_04737_),
    .B1(_03438_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_2 _10620_ (.A(_03440_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__or2_2 _10621_ (.A(_03440_),
    .B(_04764_),
    .X(_04766_));
 sky130_fd_sc_hd__mux4_2 _10622_ (.A0(_02306_),
    .A1(_02336_),
    .A2(_02291_),
    .A3(_02736_),
    .S0(_02099_),
    .S1(_04245_),
    .X(_04767_));
 sky130_fd_sc_hd__mux4_2 _10623_ (.A0(\core.cpuregs[8][15] ),
    .A1(\core.cpuregs[9][15] ),
    .A2(\core.cpuregs[10][15] ),
    .A3(\core.cpuregs[11][15] ),
    .S0(_03296_),
    .S1(_03298_),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_2 _10624_ (.A0(\core.cpuregs[14][15] ),
    .A1(\core.cpuregs[15][15] ),
    .S(_03320_),
    .X(_04769_));
 sky130_fd_sc_hd__mux2_2 _10625_ (.A0(\core.cpuregs[12][15] ),
    .A1(\core.cpuregs[13][15] ),
    .S(_03319_),
    .X(_04770_));
 sky130_fd_sc_hd__a21o_2 _10626_ (.A1(_03284_),
    .A2(_04770_),
    .B1(_03288_),
    .X(_04771_));
 sky130_fd_sc_hd__a21o_2 _10627_ (.A1(_04328_),
    .A2(_04769_),
    .B1(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__o211a_2 _10628_ (.A1(_04325_),
    .A2(_04768_),
    .B1(_04772_),
    .C1(_04508_),
    .X(_04773_));
 sky130_fd_sc_hd__mux4_2 _10629_ (.A0(\core.cpuregs[4][15] ),
    .A1(\core.cpuregs[5][15] ),
    .A2(\core.cpuregs[6][15] ),
    .A3(\core.cpuregs[7][15] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_04774_));
 sky130_fd_sc_hd__mux2_2 _10630_ (.A0(\core.cpuregs[2][15] ),
    .A1(\core.cpuregs[3][15] ),
    .S(_03329_),
    .X(_04775_));
 sky130_fd_sc_hd__mux2_2 _10631_ (.A0(\core.cpuregs[0][15] ),
    .A1(\core.cpuregs[1][15] ),
    .S(_04306_),
    .X(_04776_));
 sky130_fd_sc_hd__a21o_2 _10632_ (.A1(_04512_),
    .A2(_04776_),
    .B1(_03267_),
    .X(_04777_));
 sky130_fd_sc_hd__a21o_2 _10633_ (.A1(_03326_),
    .A2(_04775_),
    .B1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__o211a_2 _10634_ (.A1(_04259_),
    .A2(_04774_),
    .B1(_04778_),
    .C1(_04408_),
    .X(_04779_));
 sky130_fd_sc_hd__or3_2 _10635_ (.A(_04500_),
    .B(_04773_),
    .C(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__mux4_2 _10636_ (.A0(\core.cpuregs[16][15] ),
    .A1(\core.cpuregs[17][15] ),
    .A2(\core.cpuregs[18][15] ),
    .A3(\core.cpuregs[19][15] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04781_));
 sky130_fd_sc_hd__mux2_2 _10637_ (.A0(\core.cpuregs[22][15] ),
    .A1(\core.cpuregs[23][15] ),
    .S(_04592_),
    .X(_04782_));
 sky130_fd_sc_hd__mux2_2 _10638_ (.A0(\core.cpuregs[20][15] ),
    .A1(\core.cpuregs[21][15] ),
    .S(_04524_),
    .X(_04783_));
 sky130_fd_sc_hd__a21o_2 _10639_ (.A1(_04523_),
    .A2(_04783_),
    .B1(_04526_),
    .X(_04784_));
 sky130_fd_sc_hd__a21o_2 _10640_ (.A1(_04502_),
    .A2(_04782_),
    .B1(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__o211a_2 _10641_ (.A1(_04519_),
    .A2(_04781_),
    .B1(_04785_),
    .C1(_04529_),
    .X(_04786_));
 sky130_fd_sc_hd__mux4_2 _10642_ (.A0(\core.cpuregs[24][15] ),
    .A1(\core.cpuregs[25][15] ),
    .A2(\core.cpuregs[26][15] ),
    .A3(\core.cpuregs[27][15] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_04787_));
 sky130_fd_sc_hd__mux2_2 _10643_ (.A0(\core.cpuregs[30][15] ),
    .A1(\core.cpuregs[31][15] ),
    .S(_04437_),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_2 _10644_ (.A0(\core.cpuregs[28][15] ),
    .A1(\core.cpuregs[29][15] ),
    .S(_04600_),
    .X(_04789_));
 sky130_fd_sc_hd__a21o_2 _10645_ (.A1(_04403_),
    .A2(_04789_),
    .B1(_04536_),
    .X(_04790_));
 sky130_fd_sc_hd__a21o_2 _10646_ (.A1(_04533_),
    .A2(_04788_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__o211a_2 _10647_ (.A1(_04531_),
    .A2(_04787_),
    .B1(_04791_),
    .C1(_03335_),
    .X(_04792_));
 sky130_fd_sc_hd__or3_2 _10648_ (.A(_04518_),
    .B(_04786_),
    .C(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a32o_2 _10649_ (.A1(_04499_),
    .A2(_04780_),
    .A3(_04793_),
    .B1(_04541_),
    .B2(\core.reg_pc[15] ),
    .X(_04794_));
 sky130_fd_sc_hd__a22o_2 _10650_ (.A1(_02545_),
    .A2(_04767_),
    .B1(_04794_),
    .B2(_04543_),
    .X(_04795_));
 sky130_fd_sc_hd__a31o_2 _10651_ (.A1(_02235_),
    .A2(_04765_),
    .A3(_04766_),
    .B1(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__mux2_2 _10652_ (.A0(_04796_),
    .A1(_02345_),
    .S(_04639_),
    .X(_04797_));
 sky130_fd_sc_hd__buf_1 _10653_ (.A(_04797_),
    .X(_00258_));
 sky130_fd_sc_hd__nand2_2 _10654_ (.A(_03405_),
    .B(_03442_),
    .Y(_04798_));
 sky130_fd_sc_hd__nand2_2 _10655_ (.A(_03444_),
    .B(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__or2_2 _10656_ (.A(_03444_),
    .B(_04798_),
    .X(_04800_));
 sky130_fd_sc_hd__mux2_2 _10657_ (.A0(_02345_),
    .A1(_02293_),
    .S(_03469_),
    .X(_04801_));
 sky130_fd_sc_hd__mux2_2 _10658_ (.A0(_02315_),
    .A1(_02277_),
    .S(_03469_),
    .X(_04802_));
 sky130_fd_sc_hd__mux2_2 _10659_ (.A0(_04801_),
    .A1(_04802_),
    .S(_02099_),
    .X(_04803_));
 sky130_fd_sc_hd__a32o_2 _10660_ (.A1(_02041_),
    .A2(_04799_),
    .A3(_04800_),
    .B1(_04803_),
    .B2(_04244_),
    .X(_04804_));
 sky130_fd_sc_hd__mux4_2 _10661_ (.A0(\core.cpuregs[8][16] ),
    .A1(\core.cpuregs[9][16] ),
    .A2(\core.cpuregs[10][16] ),
    .A3(\core.cpuregs[11][16] ),
    .S0(_04262_),
    .S1(_04220_),
    .X(_04805_));
 sky130_fd_sc_hd__mux2_2 _10662_ (.A0(\core.cpuregs[14][16] ),
    .A1(\core.cpuregs[15][16] ),
    .S(_04385_),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_2 _10663_ (.A0(\core.cpuregs[12][16] ),
    .A1(\core.cpuregs[13][16] ),
    .S(_04326_),
    .X(_04807_));
 sky130_fd_sc_hd__a21o_2 _10664_ (.A1(_04404_),
    .A2(_04807_),
    .B1(_03332_),
    .X(_04808_));
 sky130_fd_sc_hd__a21o_2 _10665_ (.A1(_04467_),
    .A2(_04806_),
    .B1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__o211a_2 _10666_ (.A1(_04254_),
    .A2(_04805_),
    .B1(_04809_),
    .C1(_04228_),
    .X(_04810_));
 sky130_fd_sc_hd__mux4_2 _10667_ (.A0(\core.cpuregs[4][16] ),
    .A1(\core.cpuregs[5][16] ),
    .A2(\core.cpuregs[6][16] ),
    .A3(\core.cpuregs[7][16] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_2 _10668_ (.A0(\core.cpuregs[2][16] ),
    .A1(\core.cpuregs[3][16] ),
    .S(_03273_),
    .X(_04812_));
 sky130_fd_sc_hd__mux2_2 _10669_ (.A0(\core.cpuregs[0][16] ),
    .A1(\core.cpuregs[1][16] ),
    .S(_04279_),
    .X(_04813_));
 sky130_fd_sc_hd__a21o_2 _10670_ (.A1(_04469_),
    .A2(_04813_),
    .B1(_04281_),
    .X(_04814_));
 sky130_fd_sc_hd__a21o_2 _10671_ (.A1(_04285_),
    .A2(_04812_),
    .B1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__o211a_2 _10672_ (.A1(_04267_),
    .A2(_04811_),
    .B1(_04815_),
    .C1(_04240_),
    .X(_04816_));
 sky130_fd_sc_hd__or3_2 _10673_ (.A(_04265_),
    .B(_04810_),
    .C(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__mux4_2 _10674_ (.A0(\core.cpuregs[28][16] ),
    .A1(\core.cpuregs[29][16] ),
    .A2(\core.cpuregs[30][16] ),
    .A3(\core.cpuregs[31][16] ),
    .S0(_04233_),
    .S1(_04237_),
    .X(_04818_));
 sky130_fd_sc_hd__mux4_2 _10675_ (.A0(\core.cpuregs[24][16] ),
    .A1(\core.cpuregs[25][16] ),
    .A2(\core.cpuregs[26][16] ),
    .A3(\core.cpuregs[27][16] ),
    .S0(_04482_),
    .S1(_04434_),
    .X(_04819_));
 sky130_fd_sc_hd__mux4_2 _10676_ (.A0(\core.cpuregs[20][16] ),
    .A1(\core.cpuregs[21][16] ),
    .A2(\core.cpuregs[22][16] ),
    .A3(\core.cpuregs[23][16] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_04820_));
 sky130_fd_sc_hd__mux4_2 _10677_ (.A0(\core.cpuregs[16][16] ),
    .A1(\core.cpuregs[17][16] ),
    .A2(\core.cpuregs[18][16] ),
    .A3(\core.cpuregs[19][16] ),
    .S0(_04236_),
    .S1(_04400_),
    .X(_04821_));
 sky130_fd_sc_hd__mux4_2 _10678_ (.A0(_04818_),
    .A1(_04819_),
    .A2(_04820_),
    .A3(_04821_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_04822_));
 sky130_fd_sc_hd__o21a_2 _10679_ (.A1(_04242_),
    .A2(_04822_),
    .B1(_04293_),
    .X(_04823_));
 sky130_fd_sc_hd__a221o_2 _10680_ (.A1(\core.reg_pc[16] ),
    .A2(_03340_),
    .B1(_04817_),
    .B2(_04823_),
    .C1(_04491_),
    .X(_04824_));
 sky130_fd_sc_hd__o21a_2 _10681_ (.A1(_04424_),
    .A2(_04804_),
    .B1(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__mux2_2 _10682_ (.A0(_04825_),
    .A1(_02291_),
    .S(_04639_),
    .X(_04826_));
 sky130_fd_sc_hd__buf_1 _10683_ (.A(_04826_),
    .X(_00259_));
 sky130_fd_sc_hd__nand2_2 _10684_ (.A(_03372_),
    .B(_04799_),
    .Y(_04827_));
 sky130_fd_sc_hd__xor2_2 _10685_ (.A(_04827_),
    .B(_03445_),
    .X(_04828_));
 sky130_fd_sc_hd__mux4_2 _10686_ (.A0(_02312_),
    .A1(_02281_),
    .A2(_02291_),
    .A3(_02298_),
    .S0(_04298_),
    .S1(_04575_),
    .X(_04829_));
 sky130_fd_sc_hd__mux4_2 _10687_ (.A0(\core.cpuregs[8][17] ),
    .A1(\core.cpuregs[9][17] ),
    .A2(\core.cpuregs[10][17] ),
    .A3(\core.cpuregs[11][17] ),
    .S0(_04261_),
    .S1(_04219_),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_2 _10688_ (.A0(\core.cpuregs[14][17] ),
    .A1(\core.cpuregs[15][17] ),
    .S(_04307_),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_2 _10689_ (.A0(\core.cpuregs[12][17] ),
    .A1(\core.cpuregs[13][17] ),
    .S(_04317_),
    .X(_04832_));
 sky130_fd_sc_hd__a21o_2 _10690_ (.A1(_04403_),
    .A2(_04832_),
    .B1(_04536_),
    .X(_04833_));
 sky130_fd_sc_hd__a21o_2 _10691_ (.A1(_04533_),
    .A2(_04831_),
    .B1(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__o211a_2 _10692_ (.A1(_04531_),
    .A2(_04830_),
    .B1(_04834_),
    .C1(_03292_),
    .X(_04835_));
 sky130_fd_sc_hd__mux4_2 _10693_ (.A0(\core.cpuregs[4][17] ),
    .A1(\core.cpuregs[5][17] ),
    .A2(\core.cpuregs[6][17] ),
    .A3(\core.cpuregs[7][17] ),
    .S0(_04261_),
    .S1(_03278_),
    .X(_04836_));
 sky130_fd_sc_hd__mux2_2 _10694_ (.A0(\core.cpuregs[2][17] ),
    .A1(\core.cpuregs[3][17] ),
    .S(_04307_),
    .X(_04837_));
 sky130_fd_sc_hd__mux2_2 _10695_ (.A0(\core.cpuregs[0][17] ),
    .A1(\core.cpuregs[1][17] ),
    .S(_04317_),
    .X(_04838_));
 sky130_fd_sc_hd__a21o_2 _10696_ (.A1(_04276_),
    .A2(_04838_),
    .B1(_03314_),
    .X(_04839_));
 sky130_fd_sc_hd__a21o_2 _10697_ (.A1(_04387_),
    .A2(_04837_),
    .B1(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__o211a_2 _10698_ (.A1(_04266_),
    .A2(_04836_),
    .B1(_04840_),
    .C1(_03309_),
    .X(_04841_));
 sky130_fd_sc_hd__or3_2 _10699_ (.A(_03266_),
    .B(_04835_),
    .C(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__mux4_2 _10700_ (.A0(\core.cpuregs[16][17] ),
    .A1(\core.cpuregs[17][17] ),
    .A2(\core.cpuregs[18][17] ),
    .A3(\core.cpuregs[19][17] ),
    .S0(_04261_),
    .S1(_03278_),
    .X(_04843_));
 sky130_fd_sc_hd__mux2_2 _10701_ (.A0(\core.cpuregs[22][17] ),
    .A1(\core.cpuregs[23][17] ),
    .S(_04307_),
    .X(_04844_));
 sky130_fd_sc_hd__mux2_2 _10702_ (.A0(\core.cpuregs[20][17] ),
    .A1(\core.cpuregs[21][17] ),
    .S(_04317_),
    .X(_04845_));
 sky130_fd_sc_hd__a21o_2 _10703_ (.A1(_04276_),
    .A2(_04845_),
    .B1(_03289_),
    .X(_04846_));
 sky130_fd_sc_hd__a21o_2 _10704_ (.A1(_04387_),
    .A2(_04844_),
    .B1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__o211a_2 _10705_ (.A1(_03269_),
    .A2(_04843_),
    .B1(_04847_),
    .C1(_03309_),
    .X(_04848_));
 sky130_fd_sc_hd__mux4_2 _10706_ (.A0(\core.cpuregs[24][17] ),
    .A1(\core.cpuregs[25][17] ),
    .A2(\core.cpuregs[26][17] ),
    .A3(\core.cpuregs[27][17] ),
    .S0(_03281_),
    .S1(_03278_),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_2 _10707_ (.A0(\core.cpuregs[30][17] ),
    .A1(\core.cpuregs[31][17] ),
    .S(_04326_),
    .X(_04850_));
 sky130_fd_sc_hd__mux2_2 _10708_ (.A0(\core.cpuregs[28][17] ),
    .A1(\core.cpuregs[29][17] ),
    .S(_03271_),
    .X(_04851_));
 sky130_fd_sc_hd__a21o_2 _10709_ (.A1(_04276_),
    .A2(_04851_),
    .B1(_03289_),
    .X(_04852_));
 sky130_fd_sc_hd__a21o_2 _10710_ (.A1(_04387_),
    .A2(_04850_),
    .B1(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__o211a_2 _10711_ (.A1(_03269_),
    .A2(_04849_),
    .B1(_04853_),
    .C1(_03292_),
    .X(_04854_));
 sky130_fd_sc_hd__or3_2 _10712_ (.A(_03313_),
    .B(_04848_),
    .C(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a32o_2 _10713_ (.A1(_04293_),
    .A2(_04842_),
    .A3(_04855_),
    .B1(_04253_),
    .B2(\core.reg_pc[17] ),
    .X(_04856_));
 sky130_fd_sc_hd__a22o_2 _10714_ (.A1(_04244_),
    .A2(_04829_),
    .B1(_04856_),
    .B2(_03262_),
    .X(_04857_));
 sky130_fd_sc_hd__a21o_2 _10715_ (.A1(_02235_),
    .A2(_04828_),
    .B1(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__mux2_2 _10716_ (.A0(_04858_),
    .A1(_02293_),
    .S(_04639_),
    .X(_04859_));
 sky130_fd_sc_hd__buf_1 _10717_ (.A(_04859_),
    .X(_00260_));
 sky130_fd_sc_hd__a31o_2 _10718_ (.A1(_03371_),
    .A2(_03372_),
    .A3(_04799_),
    .B1(_03373_),
    .X(_04860_));
 sky130_fd_sc_hd__xor2_2 _10719_ (.A(_03377_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__mux2_2 _10720_ (.A0(_02736_),
    .A1(_02293_),
    .S(_04613_),
    .X(_04862_));
 sky130_fd_sc_hd__mux2_2 _10721_ (.A0(_02306_),
    .A1(_02408_),
    .S(_03469_),
    .X(_04863_));
 sky130_fd_sc_hd__mux2_2 _10722_ (.A0(_04862_),
    .A1(_04863_),
    .S(_03344_),
    .X(_04864_));
 sky130_fd_sc_hd__a22o_2 _10723_ (.A1(_02042_),
    .A2(_04861_),
    .B1(_04864_),
    .B2(_04377_),
    .X(_04865_));
 sky130_fd_sc_hd__mux4_2 _10724_ (.A0(\core.cpuregs[8][18] ),
    .A1(\core.cpuregs[9][18] ),
    .A2(\core.cpuregs[10][18] ),
    .A3(\core.cpuregs[11][18] ),
    .S0(_04262_),
    .S1(_04220_),
    .X(_04866_));
 sky130_fd_sc_hd__mux2_2 _10725_ (.A0(\core.cpuregs[14][18] ),
    .A1(\core.cpuregs[15][18] ),
    .S(_04385_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_2 _10726_ (.A0(\core.cpuregs[12][18] ),
    .A1(\core.cpuregs[13][18] ),
    .S(_04326_),
    .X(_04868_));
 sky130_fd_sc_hd__a21o_2 _10727_ (.A1(_04404_),
    .A2(_04868_),
    .B1(_03332_),
    .X(_04869_));
 sky130_fd_sc_hd__a21o_2 _10728_ (.A1(_03327_),
    .A2(_04867_),
    .B1(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__o211a_2 _10729_ (.A1(_04254_),
    .A2(_04866_),
    .B1(_04870_),
    .C1(_03336_),
    .X(_04871_));
 sky130_fd_sc_hd__mux4_2 _10730_ (.A0(\core.cpuregs[4][18] ),
    .A1(\core.cpuregs[5][18] ),
    .A2(\core.cpuregs[6][18] ),
    .A3(\core.cpuregs[7][18] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_04872_));
 sky130_fd_sc_hd__mux2_2 _10731_ (.A0(\core.cpuregs[2][18] ),
    .A1(\core.cpuregs[3][18] ),
    .S(_04446_),
    .X(_04873_));
 sky130_fd_sc_hd__mux2_2 _10732_ (.A0(\core.cpuregs[0][18] ),
    .A1(\core.cpuregs[1][18] ),
    .S(_04279_),
    .X(_04874_));
 sky130_fd_sc_hd__a21o_2 _10733_ (.A1(_04469_),
    .A2(_04874_),
    .B1(_04281_),
    .X(_04875_));
 sky130_fd_sc_hd__a21o_2 _10734_ (.A1(_04285_),
    .A2(_04873_),
    .B1(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__o211a_2 _10735_ (.A1(_04260_),
    .A2(_04872_),
    .B1(_04876_),
    .C1(_04487_),
    .X(_04877_));
 sky130_fd_sc_hd__or3_2 _10736_ (.A(_04265_),
    .B(_04871_),
    .C(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__mux4_2 _10737_ (.A0(\core.cpuregs[28][18] ),
    .A1(\core.cpuregs[29][18] ),
    .A2(\core.cpuregs[30][18] ),
    .A3(\core.cpuregs[31][18] ),
    .S0(_04233_),
    .S1(_04237_),
    .X(_04879_));
 sky130_fd_sc_hd__mux4_2 _10738_ (.A0(\core.cpuregs[24][18] ),
    .A1(\core.cpuregs[25][18] ),
    .A2(\core.cpuregs[26][18] ),
    .A3(\core.cpuregs[27][18] ),
    .S0(_04482_),
    .S1(_03299_),
    .X(_04880_));
 sky130_fd_sc_hd__mux4_2 _10739_ (.A0(\core.cpuregs[20][18] ),
    .A1(\core.cpuregs[21][18] ),
    .A2(\core.cpuregs[22][18] ),
    .A3(\core.cpuregs[23][18] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_04881_));
 sky130_fd_sc_hd__mux4_2 _10740_ (.A0(\core.cpuregs[16][18] ),
    .A1(\core.cpuregs[17][18] ),
    .A2(\core.cpuregs[18][18] ),
    .A3(\core.cpuregs[19][18] ),
    .S0(_04236_),
    .S1(_04400_),
    .X(_04882_));
 sky130_fd_sc_hd__mux4_2 _10741_ (.A0(_04879_),
    .A1(_04880_),
    .A2(_04881_),
    .A3(_04882_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_04883_));
 sky130_fd_sc_hd__o21a_2 _10742_ (.A1(_04242_),
    .A2(_04883_),
    .B1(_04293_),
    .X(_04884_));
 sky130_fd_sc_hd__a221o_2 _10743_ (.A1(\core.reg_pc[18] ),
    .A2(_04253_),
    .B1(_04878_),
    .B2(_04884_),
    .C1(_04491_),
    .X(_04885_));
 sky130_fd_sc_hd__o21a_2 _10744_ (.A1(_04424_),
    .A2(_04865_),
    .B1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__mux2_2 _10745_ (.A0(_04886_),
    .A1(_02298_),
    .S(_04639_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_1 _10746_ (.A(_04887_),
    .X(_00261_));
 sky130_fd_sc_hd__o21a_2 _10747_ (.A1(_03377_),
    .A2(_04860_),
    .B1(_03370_),
    .X(_04888_));
 sky130_fd_sc_hd__or3_2 _10748_ (.A(_03375_),
    .B(_03369_),
    .C(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__o21ai_2 _10749_ (.A1(_03375_),
    .A2(_03369_),
    .B1(_04888_),
    .Y(_04890_));
 sky130_fd_sc_hd__mux4_2 _10750_ (.A0(_02345_),
    .A1(_02270_),
    .A2(_02298_),
    .A3(_02277_),
    .S0(_04298_),
    .S1(_04575_),
    .X(_04891_));
 sky130_fd_sc_hd__mux4_2 _10751_ (.A0(\core.cpuregs[8][19] ),
    .A1(\core.cpuregs[9][19] ),
    .A2(\core.cpuregs[10][19] ),
    .A3(\core.cpuregs[11][19] ),
    .S0(_03296_),
    .S1(_03298_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_2 _10752_ (.A0(\core.cpuregs[14][19] ),
    .A1(\core.cpuregs[15][19] ),
    .S(_03320_),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_2 _10753_ (.A0(\core.cpuregs[12][19] ),
    .A1(\core.cpuregs[13][19] ),
    .S(_03319_),
    .X(_04894_));
 sky130_fd_sc_hd__a21o_2 _10754_ (.A1(_03284_),
    .A2(_04894_),
    .B1(_03288_),
    .X(_04895_));
 sky130_fd_sc_hd__a21o_2 _10755_ (.A1(_04328_),
    .A2(_04893_),
    .B1(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__o211a_2 _10756_ (.A1(_04325_),
    .A2(_04892_),
    .B1(_04896_),
    .C1(_04508_),
    .X(_04897_));
 sky130_fd_sc_hd__mux4_2 _10757_ (.A0(\core.cpuregs[4][19] ),
    .A1(\core.cpuregs[5][19] ),
    .A2(\core.cpuregs[6][19] ),
    .A3(\core.cpuregs[7][19] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_04898_));
 sky130_fd_sc_hd__mux2_2 _10758_ (.A0(\core.cpuregs[2][19] ),
    .A1(\core.cpuregs[3][19] ),
    .S(_03304_),
    .X(_04899_));
 sky130_fd_sc_hd__mux2_2 _10759_ (.A0(\core.cpuregs[0][19] ),
    .A1(\core.cpuregs[1][19] ),
    .S(_04306_),
    .X(_04900_));
 sky130_fd_sc_hd__a21o_2 _10760_ (.A1(_04512_),
    .A2(_04900_),
    .B1(_03267_),
    .X(_04901_));
 sky130_fd_sc_hd__a21o_2 _10761_ (.A1(_04521_),
    .A2(_04899_),
    .B1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__o211a_2 _10762_ (.A1(_04259_),
    .A2(_04898_),
    .B1(_04902_),
    .C1(_04408_),
    .X(_04903_));
 sky130_fd_sc_hd__or3_2 _10763_ (.A(_04500_),
    .B(_04897_),
    .C(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__mux4_2 _10764_ (.A0(\core.cpuregs[16][19] ),
    .A1(\core.cpuregs[17][19] ),
    .A2(\core.cpuregs[18][19] ),
    .A3(\core.cpuregs[19][19] ),
    .S0(_04314_),
    .S1(_04315_),
    .X(_04905_));
 sky130_fd_sc_hd__mux2_2 _10765_ (.A0(\core.cpuregs[22][19] ),
    .A1(\core.cpuregs[23][19] ),
    .S(_04592_),
    .X(_04906_));
 sky130_fd_sc_hd__mux2_2 _10766_ (.A0(\core.cpuregs[20][19] ),
    .A1(\core.cpuregs[21][19] ),
    .S(_04524_),
    .X(_04907_));
 sky130_fd_sc_hd__a21o_2 _10767_ (.A1(_04504_),
    .A2(_04907_),
    .B1(_04526_),
    .X(_04908_));
 sky130_fd_sc_hd__a21o_2 _10768_ (.A1(_04502_),
    .A2(_04906_),
    .B1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__o211a_2 _10769_ (.A1(_04519_),
    .A2(_04905_),
    .B1(_04909_),
    .C1(_04529_),
    .X(_04910_));
 sky130_fd_sc_hd__mux4_2 _10770_ (.A0(\core.cpuregs[24][19] ),
    .A1(\core.cpuregs[25][19] ),
    .A2(\core.cpuregs[26][19] ),
    .A3(\core.cpuregs[27][19] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_04911_));
 sky130_fd_sc_hd__mux2_2 _10771_ (.A0(\core.cpuregs[30][19] ),
    .A1(\core.cpuregs[31][19] ),
    .S(_04437_),
    .X(_04912_));
 sky130_fd_sc_hd__mux2_2 _10772_ (.A0(\core.cpuregs[28][19] ),
    .A1(\core.cpuregs[29][19] ),
    .S(_04600_),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_2 _10773_ (.A1(_04403_),
    .A2(_04913_),
    .B1(_04536_),
    .X(_04914_));
 sky130_fd_sc_hd__a21o_2 _10774_ (.A1(_04533_),
    .A2(_04912_),
    .B1(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__o211a_2 _10775_ (.A1(_04531_),
    .A2(_04911_),
    .B1(_04915_),
    .C1(_03335_),
    .X(_04916_));
 sky130_fd_sc_hd__or3_2 _10776_ (.A(_04518_),
    .B(_04910_),
    .C(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__a32o_2 _10777_ (.A1(_04499_),
    .A2(_04904_),
    .A3(_04917_),
    .B1(_04541_),
    .B2(\core.reg_pc[19] ),
    .X(_04918_));
 sky130_fd_sc_hd__a22o_2 _10778_ (.A1(_02545_),
    .A2(_04891_),
    .B1(_04918_),
    .B2(_04543_),
    .X(_04919_));
 sky130_fd_sc_hd__a31o_2 _10779_ (.A1(_02235_),
    .A2(_04889_),
    .A3(_04890_),
    .B1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__mux2_2 _10780_ (.A0(_04920_),
    .A1(_02736_),
    .S(_04639_),
    .X(_04921_));
 sky130_fd_sc_hd__buf_1 _10781_ (.A(_04921_),
    .X(_00262_));
 sky130_fd_sc_hd__o21a_2 _10782_ (.A1(_03369_),
    .A2(_04888_),
    .B1(_03379_),
    .X(_04922_));
 sky130_fd_sc_hd__nand2_2 _10783_ (.A(_03365_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__o21a_2 _10784_ (.A1(_03365_),
    .A2(_04922_),
    .B1(_02041_),
    .X(_04924_));
 sky130_fd_sc_hd__mux4_2 _10785_ (.A0(_02256_),
    .A1(_02281_),
    .A2(_02291_),
    .A3(_02736_),
    .S0(_04575_),
    .S1(_03343_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_2 _10786_ (.A1(_04923_),
    .A2(_04924_),
    .B1(_04925_),
    .B2(_04377_),
    .X(_04926_));
 sky130_fd_sc_hd__mux4_2 _10787_ (.A0(\core.cpuregs[8][20] ),
    .A1(\core.cpuregs[9][20] ),
    .A2(\core.cpuregs[10][20] ),
    .A3(\core.cpuregs[11][20] ),
    .S0(_04262_),
    .S1(_04220_),
    .X(_04927_));
 sky130_fd_sc_hd__mux2_2 _10788_ (.A0(\core.cpuregs[14][20] ),
    .A1(\core.cpuregs[15][20] ),
    .S(_04385_),
    .X(_04928_));
 sky130_fd_sc_hd__mux2_2 _10789_ (.A0(\core.cpuregs[12][20] ),
    .A1(\core.cpuregs[13][20] ),
    .S(_04326_),
    .X(_04929_));
 sky130_fd_sc_hd__a21o_2 _10790_ (.A1(_04404_),
    .A2(_04929_),
    .B1(_03332_),
    .X(_04930_));
 sky130_fd_sc_hd__a21o_2 _10791_ (.A1(_03327_),
    .A2(_04928_),
    .B1(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__o211a_2 _10792_ (.A1(_04254_),
    .A2(_04927_),
    .B1(_04931_),
    .C1(_03336_),
    .X(_04932_));
 sky130_fd_sc_hd__mux4_2 _10793_ (.A0(\core.cpuregs[4][20] ),
    .A1(\core.cpuregs[5][20] ),
    .A2(\core.cpuregs[6][20] ),
    .A3(\core.cpuregs[7][20] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_2 _10794_ (.A0(\core.cpuregs[2][20] ),
    .A1(\core.cpuregs[3][20] ),
    .S(_04446_),
    .X(_04934_));
 sky130_fd_sc_hd__mux2_2 _10795_ (.A0(\core.cpuregs[0][20] ),
    .A1(\core.cpuregs[1][20] ),
    .S(_04279_),
    .X(_04935_));
 sky130_fd_sc_hd__a21o_2 _10796_ (.A1(_04469_),
    .A2(_04935_),
    .B1(_04281_),
    .X(_04936_));
 sky130_fd_sc_hd__a21o_2 _10797_ (.A1(_04285_),
    .A2(_04934_),
    .B1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__o211a_2 _10798_ (.A1(_04260_),
    .A2(_04933_),
    .B1(_04937_),
    .C1(_04487_),
    .X(_04938_));
 sky130_fd_sc_hd__or3_2 _10799_ (.A(_04265_),
    .B(_04932_),
    .C(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__mux4_2 _10800_ (.A0(\core.cpuregs[28][20] ),
    .A1(\core.cpuregs[29][20] ),
    .A2(\core.cpuregs[30][20] ),
    .A3(\core.cpuregs[31][20] ),
    .S0(_04233_),
    .S1(_04237_),
    .X(_04940_));
 sky130_fd_sc_hd__mux4_2 _10801_ (.A0(\core.cpuregs[24][20] ),
    .A1(\core.cpuregs[25][20] ),
    .A2(\core.cpuregs[26][20] ),
    .A3(\core.cpuregs[27][20] ),
    .S0(_04482_),
    .S1(_03299_),
    .X(_04941_));
 sky130_fd_sc_hd__mux4_2 _10802_ (.A0(\core.cpuregs[20][20] ),
    .A1(\core.cpuregs[21][20] ),
    .A2(\core.cpuregs[22][20] ),
    .A3(\core.cpuregs[23][20] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_04942_));
 sky130_fd_sc_hd__mux4_2 _10803_ (.A0(\core.cpuregs[16][20] ),
    .A1(\core.cpuregs[17][20] ),
    .A2(\core.cpuregs[18][20] ),
    .A3(\core.cpuregs[19][20] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_04943_));
 sky130_fd_sc_hd__mux4_2 _10804_ (.A0(_04940_),
    .A1(_04941_),
    .A2(_04942_),
    .A3(_04943_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_04944_));
 sky130_fd_sc_hd__o21a_2 _10805_ (.A1(_04242_),
    .A2(_04944_),
    .B1(_04293_),
    .X(_04945_));
 sky130_fd_sc_hd__a221o_2 _10806_ (.A1(\core.reg_pc[20] ),
    .A2(_04253_),
    .B1(_04939_),
    .B2(_04945_),
    .C1(_04491_),
    .X(_04946_));
 sky130_fd_sc_hd__o21a_2 _10807_ (.A1(_04424_),
    .A2(_04926_),
    .B1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__buf_1 _10808_ (.A(_03473_),
    .X(_04948_));
 sky130_fd_sc_hd__mux2_2 _10809_ (.A0(_04947_),
    .A1(_02277_),
    .S(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__buf_1 _10810_ (.A(_04949_),
    .X(_00263_));
 sky130_fd_sc_hd__mux4_2 _10811_ (.A0(_02814_),
    .A1(_02408_),
    .A2(_02293_),
    .A3(_02277_),
    .S0(_02179_),
    .S1(_03343_),
    .X(_04950_));
 sky130_fd_sc_hd__o21a_2 _10812_ (.A1(_03365_),
    .A2(_04922_),
    .B1(_03359_),
    .X(_04951_));
 sky130_fd_sc_hd__xnor2_2 _10813_ (.A(_04951_),
    .B(_03367_),
    .Y(_04952_));
 sky130_fd_sc_hd__mux4_2 _10814_ (.A0(\core.cpuregs[8][21] ),
    .A1(\core.cpuregs[9][21] ),
    .A2(\core.cpuregs[10][21] ),
    .A3(\core.cpuregs[11][21] ),
    .S0(_03296_),
    .S1(_03274_),
    .X(_04953_));
 sky130_fd_sc_hd__mux2_2 _10815_ (.A0(\core.cpuregs[14][21] ),
    .A1(\core.cpuregs[15][21] ),
    .S(_03280_),
    .X(_04954_));
 sky130_fd_sc_hd__mux2_2 _10816_ (.A0(\core.cpuregs[12][21] ),
    .A1(\core.cpuregs[13][21] ),
    .S(_03319_),
    .X(_04955_));
 sky130_fd_sc_hd__a21o_2 _10817_ (.A1(_03284_),
    .A2(_04955_),
    .B1(_03288_),
    .X(_04956_));
 sky130_fd_sc_hd__a21o_2 _10818_ (.A1(_04328_),
    .A2(_04954_),
    .B1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__o211a_2 _10819_ (.A1(_04325_),
    .A2(_04953_),
    .B1(_04957_),
    .C1(_00008_),
    .X(_04958_));
 sky130_fd_sc_hd__mux4_2 _10820_ (.A0(\core.cpuregs[4][21] ),
    .A1(\core.cpuregs[5][21] ),
    .A2(\core.cpuregs[6][21] ),
    .A3(\core.cpuregs[7][21] ),
    .S0(_04314_),
    .S1(_04583_),
    .X(_04959_));
 sky130_fd_sc_hd__mux2_2 _10821_ (.A0(\core.cpuregs[2][21] ),
    .A1(\core.cpuregs[3][21] ),
    .S(_03304_),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_2 _10822_ (.A0(\core.cpuregs[0][21] ),
    .A1(\core.cpuregs[1][21] ),
    .S(_04524_),
    .X(_04961_));
 sky130_fd_sc_hd__a21o_2 _10823_ (.A1(_04523_),
    .A2(_04961_),
    .B1(_03267_),
    .X(_04962_));
 sky130_fd_sc_hd__a21o_2 _10824_ (.A1(_04521_),
    .A2(_04960_),
    .B1(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__o211a_2 _10825_ (.A1(_03294_),
    .A2(_04959_),
    .B1(_04963_),
    .C1(_04529_),
    .X(_04964_));
 sky130_fd_sc_hd__or3_2 _10826_ (.A(_00009_),
    .B(_04958_),
    .C(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__mux4_2 _10827_ (.A0(\core.cpuregs[16][21] ),
    .A1(\core.cpuregs[17][21] ),
    .A2(\core.cpuregs[18][21] ),
    .A3(\core.cpuregs[19][21] ),
    .S0(_04431_),
    .S1(_03298_),
    .X(_04966_));
 sky130_fd_sc_hd__mux2_2 _10828_ (.A0(\core.cpuregs[22][21] ),
    .A1(\core.cpuregs[23][21] ),
    .S(_04592_),
    .X(_04967_));
 sky130_fd_sc_hd__mux2_2 _10829_ (.A0(\core.cpuregs[20][21] ),
    .A1(\core.cpuregs[21][21] ),
    .S(_03303_),
    .X(_04968_));
 sky130_fd_sc_hd__a21o_2 _10830_ (.A1(_04504_),
    .A2(_04968_),
    .B1(_03331_),
    .X(_04969_));
 sky130_fd_sc_hd__a21o_2 _10831_ (.A1(_04502_),
    .A2(_04967_),
    .B1(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__o211a_2 _10832_ (.A1(_03315_),
    .A2(_04966_),
    .B1(_04970_),
    .C1(_03308_),
    .X(_04971_));
 sky130_fd_sc_hd__mux4_2 _10833_ (.A0(\core.cpuregs[24][21] ),
    .A1(\core.cpuregs[25][21] ),
    .A2(\core.cpuregs[26][21] ),
    .A3(\core.cpuregs[27][21] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_2 _10834_ (.A0(\core.cpuregs[30][21] ),
    .A1(\core.cpuregs[31][21] ),
    .S(_03329_),
    .X(_04973_));
 sky130_fd_sc_hd__mux2_2 _10835_ (.A0(\core.cpuregs[28][21] ),
    .A1(\core.cpuregs[29][21] ),
    .S(_04600_),
    .X(_04974_));
 sky130_fd_sc_hd__a21o_2 _10836_ (.A1(_04512_),
    .A2(_04974_),
    .B1(_04526_),
    .X(_04975_));
 sky130_fd_sc_hd__a21o_2 _10837_ (.A1(_03326_),
    .A2(_04973_),
    .B1(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__o211a_2 _10838_ (.A1(_04519_),
    .A2(_04972_),
    .B1(_04976_),
    .C1(_03335_),
    .X(_04977_));
 sky130_fd_sc_hd__or3_2 _10839_ (.A(_03312_),
    .B(_04971_),
    .C(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__a32o_2 _10840_ (.A1(_03264_),
    .A2(_04965_),
    .A3(_04978_),
    .B1(_04253_),
    .B2(\core.reg_pc[21] ),
    .X(_04979_));
 sky130_fd_sc_hd__a2bb2o_2 _10841_ (.A1_N(_02121_),
    .A2_N(_04952_),
    .B1(_04979_),
    .B2(_04543_),
    .X(_04980_));
 sky130_fd_sc_hd__a21o_2 _10842_ (.A1(_02116_),
    .A2(_04950_),
    .B1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__mux2_2 _10843_ (.A0(_04981_),
    .A1(_02281_),
    .S(_04948_),
    .X(_04982_));
 sky130_fd_sc_hd__buf_1 _10844_ (.A(_04982_),
    .X(_00264_));
 sky130_fd_sc_hd__or2_2 _10845_ (.A(_03360_),
    .B(_04951_),
    .X(_04983_));
 sky130_fd_sc_hd__a21oi_2 _10846_ (.A1(_03358_),
    .A2(_04983_),
    .B1(_03357_),
    .Y(_04984_));
 sky130_fd_sc_hd__and3_2 _10847_ (.A(_03357_),
    .B(_03358_),
    .C(_04983_),
    .X(_04985_));
 sky130_fd_sc_hd__nor3_2 _10848_ (.A(_02121_),
    .B(_04984_),
    .C(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__mux2_2 _10849_ (.A0(_02270_),
    .A1(_02281_),
    .S(_03343_),
    .X(_04987_));
 sky130_fd_sc_hd__mux2_2 _10850_ (.A0(_02422_),
    .A1(_02298_),
    .S(_04613_),
    .X(_04988_));
 sky130_fd_sc_hd__or2_2 _10851_ (.A(_04575_),
    .B(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__o211a_2 _10852_ (.A1(_03344_),
    .A2(_04987_),
    .B1(_04989_),
    .C1(_02545_),
    .X(_04990_));
 sky130_fd_sc_hd__mux4_2 _10853_ (.A0(\core.cpuregs[8][22] ),
    .A1(\core.cpuregs[9][22] ),
    .A2(\core.cpuregs[10][22] ),
    .A3(\core.cpuregs[11][22] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_2 _10854_ (.A0(\core.cpuregs[14][22] ),
    .A1(\core.cpuregs[15][22] ),
    .S(_04385_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_2 _10855_ (.A0(\core.cpuregs[12][22] ),
    .A1(\core.cpuregs[13][22] ),
    .S(_04326_),
    .X(_04993_));
 sky130_fd_sc_hd__a21o_2 _10856_ (.A1(_04404_),
    .A2(_04993_),
    .B1(_03332_),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_2 _10857_ (.A1(_03327_),
    .A2(_04992_),
    .B1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__o211a_2 _10858_ (.A1(_03316_),
    .A2(_04991_),
    .B1(_04995_),
    .C1(_03336_),
    .X(_04996_));
 sky130_fd_sc_hd__mux4_2 _10859_ (.A0(\core.cpuregs[4][22] ),
    .A1(\core.cpuregs[5][22] ),
    .A2(\core.cpuregs[6][22] ),
    .A3(\core.cpuregs[7][22] ),
    .S0(_04255_),
    .S1(_04256_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_2 _10860_ (.A0(\core.cpuregs[2][22] ),
    .A1(\core.cpuregs[3][22] ),
    .S(_04446_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_2 _10861_ (.A0(\core.cpuregs[0][22] ),
    .A1(\core.cpuregs[1][22] ),
    .S(_03272_),
    .X(_04999_));
 sky130_fd_sc_hd__a21o_2 _10862_ (.A1(_04469_),
    .A2(_04999_),
    .B1(_03268_),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_2 _10863_ (.A1(_04467_),
    .A2(_04998_),
    .B1(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__o211a_2 _10864_ (.A1(_04260_),
    .A2(_04997_),
    .B1(_05001_),
    .C1(_04487_),
    .X(_05002_));
 sky130_fd_sc_hd__or3_2 _10865_ (.A(_03266_),
    .B(_04996_),
    .C(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__mux4_2 _10866_ (.A0(\core.cpuregs[28][22] ),
    .A1(\core.cpuregs[29][22] ),
    .A2(\core.cpuregs[30][22] ),
    .A3(\core.cpuregs[31][22] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_2 _10867_ (.A0(\core.cpuregs[24][22] ),
    .A1(\core.cpuregs[25][22] ),
    .A2(\core.cpuregs[26][22] ),
    .A3(\core.cpuregs[27][22] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_05005_));
 sky130_fd_sc_hd__mux4_2 _10868_ (.A0(\core.cpuregs[20][22] ),
    .A1(\core.cpuregs[21][22] ),
    .A2(\core.cpuregs[22][22] ),
    .A3(\core.cpuregs[23][22] ),
    .S0(_04432_),
    .S1(_04434_),
    .X(_05006_));
 sky130_fd_sc_hd__mux4_2 _10869_ (.A0(\core.cpuregs[16][22] ),
    .A1(\core.cpuregs[17][22] ),
    .A2(\core.cpuregs[18][22] ),
    .A3(\core.cpuregs[19][22] ),
    .S0(_04399_),
    .S1(_04484_),
    .X(_05007_));
 sky130_fd_sc_hd__mux4_2 _10870_ (.A0(_05004_),
    .A1(_05005_),
    .A2(_05006_),
    .A3(_05007_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_05008_));
 sky130_fd_sc_hd__o21a_2 _10871_ (.A1(_03313_),
    .A2(_05008_),
    .B1(_04293_),
    .X(_05009_));
 sky130_fd_sc_hd__a221o_2 _10872_ (.A1(\core.reg_pc[22] ),
    .A2(_04253_),
    .B1(_05003_),
    .B2(_05009_),
    .C1(_04490_),
    .X(_05010_));
 sky130_fd_sc_hd__o31a_2 _10873_ (.A1(_03262_),
    .A2(_04986_),
    .A3(_04990_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_2 _10874_ (.A0(_05011_),
    .A1(_02408_),
    .S(_04948_),
    .X(_05012_));
 sky130_fd_sc_hd__buf_1 _10875_ (.A(_05012_),
    .X(_00265_));
 sky130_fd_sc_hd__a21o_2 _10876_ (.A1(_02408_),
    .A2(\core.decoded_imm[22] ),
    .B1(_04984_),
    .X(_05013_));
 sky130_fd_sc_hd__or2b_2 _10877_ (.A(_03363_),
    .B_N(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__or2b_2 _10878_ (.A(_05013_),
    .B_N(_03363_),
    .X(_05015_));
 sky130_fd_sc_hd__mux4_2 _10879_ (.A0(_02838_),
    .A1(_02256_),
    .A2(_02736_),
    .A3(_02408_),
    .S0(_02178_),
    .S1(_03343_),
    .X(_05016_));
 sky130_fd_sc_hd__mux4_2 _10880_ (.A0(\core.cpuregs[8][23] ),
    .A1(\core.cpuregs[9][23] ),
    .A2(\core.cpuregs[10][23] ),
    .A3(\core.cpuregs[11][23] ),
    .S0(_03296_),
    .S1(_03298_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_2 _10881_ (.A0(\core.cpuregs[14][23] ),
    .A1(\core.cpuregs[15][23] ),
    .S(_03320_),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_2 _10882_ (.A0(\core.cpuregs[12][23] ),
    .A1(\core.cpuregs[13][23] ),
    .S(_03319_),
    .X(_05019_));
 sky130_fd_sc_hd__a21o_2 _10883_ (.A1(_03284_),
    .A2(_05019_),
    .B1(_03288_),
    .X(_05020_));
 sky130_fd_sc_hd__a21o_2 _10884_ (.A1(_04328_),
    .A2(_05018_),
    .B1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__o211a_2 _10885_ (.A1(_04325_),
    .A2(_05017_),
    .B1(_05021_),
    .C1(_04508_),
    .X(_05022_));
 sky130_fd_sc_hd__mux4_2 _10886_ (.A0(\core.cpuregs[4][23] ),
    .A1(\core.cpuregs[5][23] ),
    .A2(\core.cpuregs[6][23] ),
    .A3(\core.cpuregs[7][23] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_05023_));
 sky130_fd_sc_hd__mux2_2 _10887_ (.A0(\core.cpuregs[2][23] ),
    .A1(\core.cpuregs[3][23] ),
    .S(_03304_),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_2 _10888_ (.A0(\core.cpuregs[0][23] ),
    .A1(\core.cpuregs[1][23] ),
    .S(_04306_),
    .X(_05025_));
 sky130_fd_sc_hd__a21o_2 _10889_ (.A1(_04523_),
    .A2(_05025_),
    .B1(_03267_),
    .X(_05026_));
 sky130_fd_sc_hd__a21o_2 _10890_ (.A1(_04521_),
    .A2(_05024_),
    .B1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__o211a_2 _10891_ (.A1(_04259_),
    .A2(_05023_),
    .B1(_05027_),
    .C1(_04408_),
    .X(_05028_));
 sky130_fd_sc_hd__or3_2 _10892_ (.A(_04500_),
    .B(_05022_),
    .C(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__mux4_2 _10893_ (.A0(\core.cpuregs[16][23] ),
    .A1(\core.cpuregs[17][23] ),
    .A2(\core.cpuregs[18][23] ),
    .A3(\core.cpuregs[19][23] ),
    .S0(_04431_),
    .S1(_04315_),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_2 _10894_ (.A0(\core.cpuregs[22][23] ),
    .A1(\core.cpuregs[23][23] ),
    .S(_04592_),
    .X(_05031_));
 sky130_fd_sc_hd__mux2_2 _10895_ (.A0(\core.cpuregs[20][23] ),
    .A1(\core.cpuregs[21][23] ),
    .S(_04524_),
    .X(_05032_));
 sky130_fd_sc_hd__a21o_2 _10896_ (.A1(_04504_),
    .A2(_05032_),
    .B1(_03331_),
    .X(_05033_));
 sky130_fd_sc_hd__a21o_2 _10897_ (.A1(_04502_),
    .A2(_05031_),
    .B1(_05033_),
    .X(_05034_));
 sky130_fd_sc_hd__o211a_2 _10898_ (.A1(_04519_),
    .A2(_05030_),
    .B1(_05034_),
    .C1(_04529_),
    .X(_05035_));
 sky130_fd_sc_hd__mux4_2 _10899_ (.A0(\core.cpuregs[24][23] ),
    .A1(\core.cpuregs[25][23] ),
    .A2(\core.cpuregs[26][23] ),
    .A3(\core.cpuregs[27][23] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_2 _10900_ (.A0(\core.cpuregs[30][23] ),
    .A1(\core.cpuregs[31][23] ),
    .S(_04437_),
    .X(_05037_));
 sky130_fd_sc_hd__mux2_2 _10901_ (.A0(\core.cpuregs[28][23] ),
    .A1(\core.cpuregs[29][23] ),
    .S(_04600_),
    .X(_05038_));
 sky130_fd_sc_hd__a21o_2 _10902_ (.A1(_04403_),
    .A2(_05038_),
    .B1(_04536_),
    .X(_05039_));
 sky130_fd_sc_hd__a21o_2 _10903_ (.A1(_04533_),
    .A2(_05037_),
    .B1(_05039_),
    .X(_05040_));
 sky130_fd_sc_hd__o211a_2 _10904_ (.A1(_04531_),
    .A2(_05036_),
    .B1(_05040_),
    .C1(_03335_),
    .X(_05041_));
 sky130_fd_sc_hd__or3_2 _10905_ (.A(_04518_),
    .B(_05035_),
    .C(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a32o_2 _10906_ (.A1(_04499_),
    .A2(_05029_),
    .A3(_05042_),
    .B1(_04541_),
    .B2(\core.reg_pc[23] ),
    .X(_05043_));
 sky130_fd_sc_hd__a22o_2 _10907_ (.A1(_02545_),
    .A2(_05016_),
    .B1(_05043_),
    .B2(_04543_),
    .X(_05044_));
 sky130_fd_sc_hd__a31o_2 _10908_ (.A1(_02235_),
    .A2(_05014_),
    .A3(_05015_),
    .B1(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__mux2_2 _10909_ (.A0(_05045_),
    .A1(_02270_),
    .S(_04948_),
    .X(_05046_));
 sky130_fd_sc_hd__buf_1 _10910_ (.A(_05046_),
    .X(_00266_));
 sky130_fd_sc_hd__xor2_2 _10911_ (.A(_03448_),
    .B(_03451_),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_2 _10912_ (.A0(_02814_),
    .A1(_02270_),
    .S(_04613_),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_2 _10913_ (.A0(_02246_),
    .A1(_02277_),
    .S(_04613_),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_2 _10914_ (.A0(_05048_),
    .A1(_05049_),
    .S(_03344_),
    .X(_05050_));
 sky130_fd_sc_hd__a22o_2 _10915_ (.A1(_02042_),
    .A2(_05047_),
    .B1(_05050_),
    .B2(_04377_),
    .X(_05051_));
 sky130_fd_sc_hd__mux4_2 _10916_ (.A0(\core.cpuregs[8][24] ),
    .A1(\core.cpuregs[9][24] ),
    .A2(\core.cpuregs[10][24] ),
    .A3(\core.cpuregs[11][24] ),
    .S0(_04262_),
    .S1(_04220_),
    .X(_05052_));
 sky130_fd_sc_hd__mux2_2 _10917_ (.A0(\core.cpuregs[14][24] ),
    .A1(\core.cpuregs[15][24] ),
    .S(_04385_),
    .X(_05053_));
 sky130_fd_sc_hd__mux2_2 _10918_ (.A0(\core.cpuregs[12][24] ),
    .A1(\core.cpuregs[13][24] ),
    .S(_04326_),
    .X(_05054_));
 sky130_fd_sc_hd__a21o_2 _10919_ (.A1(_04404_),
    .A2(_05054_),
    .B1(_03332_),
    .X(_05055_));
 sky130_fd_sc_hd__a21o_2 _10920_ (.A1(_03327_),
    .A2(_05053_),
    .B1(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__o211a_2 _10921_ (.A1(_03316_),
    .A2(_05052_),
    .B1(_05056_),
    .C1(_03336_),
    .X(_05057_));
 sky130_fd_sc_hd__mux4_2 _10922_ (.A0(\core.cpuregs[4][24] ),
    .A1(\core.cpuregs[5][24] ),
    .A2(\core.cpuregs[6][24] ),
    .A3(\core.cpuregs[7][24] ),
    .S0(_04255_),
    .S1(_04274_),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_2 _10923_ (.A0(\core.cpuregs[2][24] ),
    .A1(\core.cpuregs[3][24] ),
    .S(_04446_),
    .X(_05059_));
 sky130_fd_sc_hd__mux2_2 _10924_ (.A0(\core.cpuregs[0][24] ),
    .A1(\core.cpuregs[1][24] ),
    .S(_04279_),
    .X(_05060_));
 sky130_fd_sc_hd__a21o_2 _10925_ (.A1(_04469_),
    .A2(_05060_),
    .B1(_04281_),
    .X(_05061_));
 sky130_fd_sc_hd__a21o_2 _10926_ (.A1(_04467_),
    .A2(_05059_),
    .B1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__o211a_2 _10927_ (.A1(_04260_),
    .A2(_05058_),
    .B1(_05062_),
    .C1(_04487_),
    .X(_05063_));
 sky130_fd_sc_hd__or3_2 _10928_ (.A(_03266_),
    .B(_05057_),
    .C(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__mux4_2 _10929_ (.A0(\core.cpuregs[28][24] ),
    .A1(\core.cpuregs[29][24] ),
    .A2(\core.cpuregs[30][24] ),
    .A3(\core.cpuregs[31][24] ),
    .S0(_04233_),
    .S1(_04237_),
    .X(_05065_));
 sky130_fd_sc_hd__mux4_2 _10930_ (.A0(\core.cpuregs[24][24] ),
    .A1(\core.cpuregs[25][24] ),
    .A2(\core.cpuregs[26][24] ),
    .A3(\core.cpuregs[27][24] ),
    .S0(_04482_),
    .S1(_03299_),
    .X(_05066_));
 sky130_fd_sc_hd__mux4_2 _10931_ (.A0(\core.cpuregs[20][24] ),
    .A1(\core.cpuregs[21][24] ),
    .A2(\core.cpuregs[22][24] ),
    .A3(\core.cpuregs[23][24] ),
    .S0(_04432_),
    .S1(_04484_),
    .X(_05067_));
 sky130_fd_sc_hd__mux4_2 _10932_ (.A0(\core.cpuregs[16][24] ),
    .A1(\core.cpuregs[17][24] ),
    .A2(\core.cpuregs[18][24] ),
    .A3(\core.cpuregs[19][24] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_05068_));
 sky130_fd_sc_hd__mux4_2 _10933_ (.A0(_05065_),
    .A1(_05066_),
    .A2(_05067_),
    .A3(_05068_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_05069_));
 sky130_fd_sc_hd__o21a_2 _10934_ (.A1(_04242_),
    .A2(_05069_),
    .B1(_04293_),
    .X(_05070_));
 sky130_fd_sc_hd__a221o_2 _10935_ (.A1(\core.reg_pc[24] ),
    .A2(_04253_),
    .B1(_05064_),
    .B2(_05070_),
    .C1(_04491_),
    .X(_05071_));
 sky130_fd_sc_hd__o21a_2 _10936_ (.A1(_03262_),
    .A2(_05051_),
    .B1(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__mux2_2 _10937_ (.A0(_05072_),
    .A1(_02256_),
    .S(_04948_),
    .X(_05073_));
 sky130_fd_sc_hd__buf_1 _10938_ (.A(_05073_),
    .X(_00267_));
 sky130_fd_sc_hd__o21ai_2 _10939_ (.A1(_03448_),
    .A2(_03451_),
    .B1(_03449_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand3_2 _10940_ (.A(_03353_),
    .B(_03452_),
    .C(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__a21o_2 _10941_ (.A1(_03353_),
    .A2(_03452_),
    .B1(_05074_),
    .X(_05076_));
 sky130_fd_sc_hd__mux4_2 _10942_ (.A0(_02414_),
    .A1(_02422_),
    .A2(_02281_),
    .A3(_02256_),
    .S0(_02178_),
    .S1(_03343_),
    .X(_05077_));
 sky130_fd_sc_hd__mux4_2 _10943_ (.A0(\core.cpuregs[8][25] ),
    .A1(\core.cpuregs[9][25] ),
    .A2(\core.cpuregs[10][25] ),
    .A3(\core.cpuregs[11][25] ),
    .S0(_03296_),
    .S1(_03274_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_2 _10944_ (.A0(\core.cpuregs[14][25] ),
    .A1(\core.cpuregs[15][25] ),
    .S(_03320_),
    .X(_05079_));
 sky130_fd_sc_hd__mux2_2 _10945_ (.A0(\core.cpuregs[12][25] ),
    .A1(\core.cpuregs[13][25] ),
    .S(_03319_),
    .X(_05080_));
 sky130_fd_sc_hd__a21o_2 _10946_ (.A1(_03284_),
    .A2(_05080_),
    .B1(_03288_),
    .X(_05081_));
 sky130_fd_sc_hd__a21o_2 _10947_ (.A1(_04328_),
    .A2(_05079_),
    .B1(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__o211a_2 _10948_ (.A1(_04325_),
    .A2(_05078_),
    .B1(_05082_),
    .C1(_04508_),
    .X(_05083_));
 sky130_fd_sc_hd__mux4_2 _10949_ (.A0(\core.cpuregs[4][25] ),
    .A1(\core.cpuregs[5][25] ),
    .A2(\core.cpuregs[6][25] ),
    .A3(\core.cpuregs[7][25] ),
    .S0(_04235_),
    .S1(_04583_),
    .X(_05084_));
 sky130_fd_sc_hd__mux2_2 _10950_ (.A0(\core.cpuregs[2][25] ),
    .A1(\core.cpuregs[3][25] ),
    .S(_03304_),
    .X(_05085_));
 sky130_fd_sc_hd__mux2_2 _10951_ (.A0(\core.cpuregs[0][25] ),
    .A1(\core.cpuregs[1][25] ),
    .S(_04306_),
    .X(_05086_));
 sky130_fd_sc_hd__a21o_2 _10952_ (.A1(_04523_),
    .A2(_05086_),
    .B1(_03267_),
    .X(_05087_));
 sky130_fd_sc_hd__a21o_2 _10953_ (.A1(_04521_),
    .A2(_05085_),
    .B1(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__o211a_2 _10954_ (.A1(_04259_),
    .A2(_05084_),
    .B1(_05088_),
    .C1(_04408_),
    .X(_05089_));
 sky130_fd_sc_hd__or3_2 _10955_ (.A(_04500_),
    .B(_05083_),
    .C(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__mux4_2 _10956_ (.A0(\core.cpuregs[16][25] ),
    .A1(\core.cpuregs[17][25] ),
    .A2(\core.cpuregs[18][25] ),
    .A3(\core.cpuregs[19][25] ),
    .S0(_04431_),
    .S1(_04315_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_2 _10957_ (.A0(\core.cpuregs[22][25] ),
    .A1(\core.cpuregs[23][25] ),
    .S(_04592_),
    .X(_05092_));
 sky130_fd_sc_hd__mux2_2 _10958_ (.A0(\core.cpuregs[20][25] ),
    .A1(\core.cpuregs[21][25] ),
    .S(_03303_),
    .X(_05093_));
 sky130_fd_sc_hd__a21o_2 _10959_ (.A1(_04504_),
    .A2(_05093_),
    .B1(_03331_),
    .X(_05094_));
 sky130_fd_sc_hd__a21o_2 _10960_ (.A1(_04502_),
    .A2(_05092_),
    .B1(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__o211a_2 _10961_ (.A1(_03315_),
    .A2(_05091_),
    .B1(_05095_),
    .C1(_04529_),
    .X(_05096_));
 sky130_fd_sc_hd__mux4_2 _10962_ (.A0(\core.cpuregs[24][25] ),
    .A1(\core.cpuregs[25][25] ),
    .A2(\core.cpuregs[26][25] ),
    .A3(\core.cpuregs[27][25] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_05097_));
 sky130_fd_sc_hd__mux2_2 _10963_ (.A0(\core.cpuregs[30][25] ),
    .A1(\core.cpuregs[31][25] ),
    .S(_04437_),
    .X(_05098_));
 sky130_fd_sc_hd__mux2_2 _10964_ (.A0(\core.cpuregs[28][25] ),
    .A1(\core.cpuregs[29][25] ),
    .S(_04600_),
    .X(_05099_));
 sky130_fd_sc_hd__a21o_2 _10965_ (.A1(_04512_),
    .A2(_05099_),
    .B1(_04526_),
    .X(_05100_));
 sky130_fd_sc_hd__a21o_2 _10966_ (.A1(_04533_),
    .A2(_05098_),
    .B1(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__o211a_2 _10967_ (.A1(_04531_),
    .A2(_05097_),
    .B1(_05101_),
    .C1(_03335_),
    .X(_05102_));
 sky130_fd_sc_hd__or3_2 _10968_ (.A(_04518_),
    .B(_05096_),
    .C(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__a32o_2 _10969_ (.A1(_04499_),
    .A2(_05090_),
    .A3(_05103_),
    .B1(_04541_),
    .B2(\core.reg_pc[25] ),
    .X(_05104_));
 sky130_fd_sc_hd__a22o_2 _10970_ (.A1(_02545_),
    .A2(_05077_),
    .B1(_05104_),
    .B2(_04543_),
    .X(_05105_));
 sky130_fd_sc_hd__a31o_2 _10971_ (.A1(_02042_),
    .A2(_05075_),
    .A3(_05076_),
    .B1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__mux2_2 _10972_ (.A0(_05106_),
    .A1(_02814_),
    .S(_04948_),
    .X(_05107_));
 sky130_fd_sc_hd__buf_1 _10973_ (.A(_05107_),
    .X(_00268_));
 sky130_fd_sc_hd__a21oi_2 _10974_ (.A1(_03353_),
    .A2(_03453_),
    .B1(_03352_),
    .Y(_05108_));
 sky130_fd_sc_hd__nor2_2 _10975_ (.A(_03454_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__mux4_2 _10976_ (.A0(_02242_),
    .A1(_02838_),
    .A2(_02408_),
    .A3(_02814_),
    .S0(_04575_),
    .S1(_03343_),
    .X(_05110_));
 sky130_fd_sc_hd__a22o_2 _10977_ (.A1(_02042_),
    .A2(_05109_),
    .B1(_05110_),
    .B2(_04377_),
    .X(_05111_));
 sky130_fd_sc_hd__mux4_2 _10978_ (.A0(\core.cpuregs[8][26] ),
    .A1(\core.cpuregs[9][26] ),
    .A2(\core.cpuregs[10][26] ),
    .A3(\core.cpuregs[11][26] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_05112_));
 sky130_fd_sc_hd__mux2_2 _10979_ (.A0(\core.cpuregs[14][26] ),
    .A1(\core.cpuregs[15][26] ),
    .S(_04385_),
    .X(_05113_));
 sky130_fd_sc_hd__mux2_2 _10980_ (.A0(\core.cpuregs[12][26] ),
    .A1(\core.cpuregs[13][26] ),
    .S(_04326_),
    .X(_05114_));
 sky130_fd_sc_hd__a21o_2 _10981_ (.A1(_04404_),
    .A2(_05114_),
    .B1(_03332_),
    .X(_05115_));
 sky130_fd_sc_hd__a21o_2 _10982_ (.A1(_03327_),
    .A2(_05113_),
    .B1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o211a_2 _10983_ (.A1(_03316_),
    .A2(_05112_),
    .B1(_05116_),
    .C1(_03336_),
    .X(_05117_));
 sky130_fd_sc_hd__mux4_2 _10984_ (.A0(\core.cpuregs[4][26] ),
    .A1(\core.cpuregs[5][26] ),
    .A2(\core.cpuregs[6][26] ),
    .A3(\core.cpuregs[7][26] ),
    .S0(_04255_),
    .S1(_04256_),
    .X(_05118_));
 sky130_fd_sc_hd__mux2_2 _10985_ (.A0(\core.cpuregs[2][26] ),
    .A1(\core.cpuregs[3][26] ),
    .S(_04446_),
    .X(_05119_));
 sky130_fd_sc_hd__mux2_2 _10986_ (.A0(\core.cpuregs[0][26] ),
    .A1(\core.cpuregs[1][26] ),
    .S(_03272_),
    .X(_05120_));
 sky130_fd_sc_hd__a21o_2 _10987_ (.A1(_04469_),
    .A2(_05120_),
    .B1(_03268_),
    .X(_05121_));
 sky130_fd_sc_hd__a21o_2 _10988_ (.A1(_04467_),
    .A2(_05119_),
    .B1(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__o211a_2 _10989_ (.A1(_04260_),
    .A2(_05118_),
    .B1(_05122_),
    .C1(_04487_),
    .X(_05123_));
 sky130_fd_sc_hd__or3_2 _10990_ (.A(_03266_),
    .B(_05117_),
    .C(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__mux4_2 _10991_ (.A0(\core.cpuregs[28][26] ),
    .A1(\core.cpuregs[29][26] ),
    .A2(\core.cpuregs[30][26] ),
    .A3(\core.cpuregs[31][26] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_05125_));
 sky130_fd_sc_hd__mux4_2 _10992_ (.A0(\core.cpuregs[24][26] ),
    .A1(\core.cpuregs[25][26] ),
    .A2(\core.cpuregs[26][26] ),
    .A3(\core.cpuregs[27][26] ),
    .S0(_04482_),
    .S1(_03299_),
    .X(_05126_));
 sky130_fd_sc_hd__mux4_2 _10993_ (.A0(\core.cpuregs[20][26] ),
    .A1(\core.cpuregs[21][26] ),
    .A2(\core.cpuregs[22][26] ),
    .A3(\core.cpuregs[23][26] ),
    .S0(_04432_),
    .S1(_04434_),
    .X(_05127_));
 sky130_fd_sc_hd__mux4_2 _10994_ (.A0(\core.cpuregs[16][26] ),
    .A1(\core.cpuregs[17][26] ),
    .A2(\core.cpuregs[18][26] ),
    .A3(\core.cpuregs[19][26] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_05128_));
 sky130_fd_sc_hd__mux4_2 _10995_ (.A0(_05125_),
    .A1(_05126_),
    .A2(_05127_),
    .A3(_05128_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_05129_));
 sky130_fd_sc_hd__o21a_2 _10996_ (.A1(_03313_),
    .A2(_05129_),
    .B1(_04293_),
    .X(_05130_));
 sky130_fd_sc_hd__a221o_2 _10997_ (.A1(\core.reg_pc[26] ),
    .A2(_04253_),
    .B1(_05124_),
    .B2(_05130_),
    .C1(_04491_),
    .X(_05131_));
 sky130_fd_sc_hd__o21a_2 _10998_ (.A1(_03262_),
    .A2(_05111_),
    .B1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_2 _10999_ (.A0(_05132_),
    .A1(_02422_),
    .S(_04948_),
    .X(_05133_));
 sky130_fd_sc_hd__buf_1 _11000_ (.A(_05133_),
    .X(_00269_));
 sky130_fd_sc_hd__nor2_2 _11001_ (.A(_03456_),
    .B(_03351_),
    .Y(_05134_));
 sky130_fd_sc_hd__xnor2_2 _11002_ (.A(_03455_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__mux4_2 _11003_ (.A0(_02237_),
    .A1(_02246_),
    .A2(_02270_),
    .A3(_02422_),
    .S0(_02178_),
    .S1(_03343_),
    .X(_05136_));
 sky130_fd_sc_hd__mux4_2 _11004_ (.A0(\core.cpuregs[8][27] ),
    .A1(\core.cpuregs[9][27] ),
    .A2(\core.cpuregs[10][27] ),
    .A3(\core.cpuregs[11][27] ),
    .S0(_04261_),
    .S1(_04219_),
    .X(_05137_));
 sky130_fd_sc_hd__mux2_2 _11005_ (.A0(\core.cpuregs[14][27] ),
    .A1(\core.cpuregs[15][27] ),
    .S(_04307_),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_2 _11006_ (.A0(\core.cpuregs[12][27] ),
    .A1(\core.cpuregs[13][27] ),
    .S(_04317_),
    .X(_05139_));
 sky130_fd_sc_hd__a21o_2 _11007_ (.A1(_04403_),
    .A2(_05139_),
    .B1(_04536_),
    .X(_05140_));
 sky130_fd_sc_hd__a21o_2 _11008_ (.A1(_04533_),
    .A2(_05138_),
    .B1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__o211a_2 _11009_ (.A1(_04531_),
    .A2(_05137_),
    .B1(_05141_),
    .C1(_03292_),
    .X(_05142_));
 sky130_fd_sc_hd__mux4_2 _11010_ (.A0(\core.cpuregs[4][27] ),
    .A1(\core.cpuregs[5][27] ),
    .A2(\core.cpuregs[6][27] ),
    .A3(\core.cpuregs[7][27] ),
    .S0(_04261_),
    .S1(_03278_),
    .X(_05143_));
 sky130_fd_sc_hd__mux2_2 _11011_ (.A0(\core.cpuregs[2][27] ),
    .A1(\core.cpuregs[3][27] ),
    .S(_04307_),
    .X(_05144_));
 sky130_fd_sc_hd__mux2_2 _11012_ (.A0(\core.cpuregs[0][27] ),
    .A1(\core.cpuregs[1][27] ),
    .S(_04317_),
    .X(_05145_));
 sky130_fd_sc_hd__a21o_2 _11013_ (.A1(_04276_),
    .A2(_05145_),
    .B1(_03314_),
    .X(_05146_));
 sky130_fd_sc_hd__a21o_2 _11014_ (.A1(_04387_),
    .A2(_05144_),
    .B1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__o211a_2 _11015_ (.A1(_04259_),
    .A2(_05143_),
    .B1(_05147_),
    .C1(_03309_),
    .X(_05148_));
 sky130_fd_sc_hd__or3_2 _11016_ (.A(_03266_),
    .B(_05142_),
    .C(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__mux4_2 _11017_ (.A0(\core.cpuregs[16][27] ),
    .A1(\core.cpuregs[17][27] ),
    .A2(\core.cpuregs[18][27] ),
    .A3(\core.cpuregs[19][27] ),
    .S0(_04261_),
    .S1(_03278_),
    .X(_05150_));
 sky130_fd_sc_hd__mux2_2 _11018_ (.A0(\core.cpuregs[22][27] ),
    .A1(\core.cpuregs[23][27] ),
    .S(_04307_),
    .X(_05151_));
 sky130_fd_sc_hd__mux2_2 _11019_ (.A0(\core.cpuregs[20][27] ),
    .A1(\core.cpuregs[21][27] ),
    .S(_04317_),
    .X(_05152_));
 sky130_fd_sc_hd__a21o_2 _11020_ (.A1(_04276_),
    .A2(_05152_),
    .B1(_04536_),
    .X(_05153_));
 sky130_fd_sc_hd__a21o_2 _11021_ (.A1(_04387_),
    .A2(_05151_),
    .B1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__o211a_2 _11022_ (.A1(_03269_),
    .A2(_05150_),
    .B1(_05154_),
    .C1(_03309_),
    .X(_05155_));
 sky130_fd_sc_hd__mux4_2 _11023_ (.A0(\core.cpuregs[24][27] ),
    .A1(\core.cpuregs[25][27] ),
    .A2(\core.cpuregs[26][27] ),
    .A3(\core.cpuregs[27][27] ),
    .S0(_03281_),
    .S1(_03278_),
    .X(_05156_));
 sky130_fd_sc_hd__mux2_2 _11024_ (.A0(\core.cpuregs[30][27] ),
    .A1(\core.cpuregs[31][27] ),
    .S(_04326_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_2 _11025_ (.A0(\core.cpuregs[28][27] ),
    .A1(\core.cpuregs[29][27] ),
    .S(_03271_),
    .X(_05158_));
 sky130_fd_sc_hd__a21o_2 _11026_ (.A1(_04276_),
    .A2(_05158_),
    .B1(_03289_),
    .X(_05159_));
 sky130_fd_sc_hd__a21o_2 _11027_ (.A1(_04387_),
    .A2(_05157_),
    .B1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__o211a_2 _11028_ (.A1(_03269_),
    .A2(_05156_),
    .B1(_05160_),
    .C1(_03292_),
    .X(_05161_));
 sky130_fd_sc_hd__or3_2 _11029_ (.A(_04518_),
    .B(_05155_),
    .C(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__a32o_2 _11030_ (.A1(_04293_),
    .A2(_05149_),
    .A3(_05162_),
    .B1(_04253_),
    .B2(\core.reg_pc[27] ),
    .X(_05163_));
 sky130_fd_sc_hd__a22o_2 _11031_ (.A1(_04244_),
    .A2(_05136_),
    .B1(_05163_),
    .B2(_04543_),
    .X(_05164_));
 sky130_fd_sc_hd__a21o_2 _11032_ (.A1(_02235_),
    .A2(_05135_),
    .B1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_2 _11033_ (.A0(_05165_),
    .A1(_02838_),
    .S(_04948_),
    .X(_05166_));
 sky130_fd_sc_hd__buf_1 _11034_ (.A(_05166_),
    .X(_00270_));
 sky130_fd_sc_hd__or3_2 _11035_ (.A(_03458_),
    .B(_03350_),
    .C(_03457_),
    .X(_05167_));
 sky130_fd_sc_hd__o21ai_2 _11036_ (.A1(_03458_),
    .A2(_03350_),
    .B1(_03457_),
    .Y(_05168_));
 sky130_fd_sc_hd__a21oi_2 _11037_ (.A1(_02237_),
    .A2(_02059_),
    .B1(_04613_),
    .Y(_05169_));
 sky130_fd_sc_hd__o21ai_2 _11038_ (.A1(_02256_),
    .A2(_04298_),
    .B1(_02099_),
    .Y(_05170_));
 sky130_fd_sc_hd__mux2_2 _11039_ (.A0(_02414_),
    .A1(_02838_),
    .S(_04613_),
    .X(_05171_));
 sky130_fd_sc_hd__a2bb2o_2 _11040_ (.A1_N(_05169_),
    .A2_N(_05170_),
    .B1(_04575_),
    .B2(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__mux4_2 _11041_ (.A0(\core.cpuregs[8][28] ),
    .A1(\core.cpuregs[9][28] ),
    .A2(\core.cpuregs[10][28] ),
    .A3(\core.cpuregs[11][28] ),
    .S0(_03296_),
    .S1(_03274_),
    .X(_05173_));
 sky130_fd_sc_hd__mux2_2 _11042_ (.A0(\core.cpuregs[14][28] ),
    .A1(\core.cpuregs[15][28] ),
    .S(_03280_),
    .X(_05174_));
 sky130_fd_sc_hd__mux2_2 _11043_ (.A0(\core.cpuregs[12][28] ),
    .A1(\core.cpuregs[13][28] ),
    .S(_03319_),
    .X(_05175_));
 sky130_fd_sc_hd__a21o_2 _11044_ (.A1(_03284_),
    .A2(_05175_),
    .B1(_03288_),
    .X(_05176_));
 sky130_fd_sc_hd__a21o_2 _11045_ (.A1(_04328_),
    .A2(_05174_),
    .B1(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__o211a_2 _11046_ (.A1(_04325_),
    .A2(_05173_),
    .B1(_05177_),
    .C1(_04508_),
    .X(_05178_));
 sky130_fd_sc_hd__mux4_2 _11047_ (.A0(\core.cpuregs[4][28] ),
    .A1(\core.cpuregs[5][28] ),
    .A2(\core.cpuregs[6][28] ),
    .A3(\core.cpuregs[7][28] ),
    .S0(_04314_),
    .S1(_04583_),
    .X(_05179_));
 sky130_fd_sc_hd__mux2_2 _11048_ (.A0(\core.cpuregs[2][28] ),
    .A1(\core.cpuregs[3][28] ),
    .S(_03304_),
    .X(_05180_));
 sky130_fd_sc_hd__mux2_2 _11049_ (.A0(\core.cpuregs[0][28] ),
    .A1(\core.cpuregs[1][28] ),
    .S(_04524_),
    .X(_05181_));
 sky130_fd_sc_hd__a21o_2 _11050_ (.A1(_04523_),
    .A2(_05181_),
    .B1(_03267_),
    .X(_05182_));
 sky130_fd_sc_hd__a21o_2 _11051_ (.A1(_04521_),
    .A2(_05180_),
    .B1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__o211a_2 _11052_ (.A1(_03294_),
    .A2(_05179_),
    .B1(_05183_),
    .C1(_04408_),
    .X(_05184_));
 sky130_fd_sc_hd__or3_2 _11053_ (.A(_04500_),
    .B(_05178_),
    .C(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__mux4_2 _11054_ (.A0(\core.cpuregs[16][28] ),
    .A1(\core.cpuregs[17][28] ),
    .A2(\core.cpuregs[18][28] ),
    .A3(\core.cpuregs[19][28] ),
    .S0(_04431_),
    .S1(_04315_),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_2 _11055_ (.A0(\core.cpuregs[22][28] ),
    .A1(\core.cpuregs[23][28] ),
    .S(_04592_),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_2 _11056_ (.A0(\core.cpuregs[20][28] ),
    .A1(\core.cpuregs[21][28] ),
    .S(_03303_),
    .X(_05188_));
 sky130_fd_sc_hd__a21o_2 _11057_ (.A1(_04504_),
    .A2(_05188_),
    .B1(_03331_),
    .X(_05189_));
 sky130_fd_sc_hd__a21o_2 _11058_ (.A1(_04502_),
    .A2(_05187_),
    .B1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__o211a_2 _11059_ (.A1(_03315_),
    .A2(_05186_),
    .B1(_05190_),
    .C1(_03308_),
    .X(_05191_));
 sky130_fd_sc_hd__mux4_2 _11060_ (.A0(\core.cpuregs[24][28] ),
    .A1(\core.cpuregs[25][28] ),
    .A2(\core.cpuregs[26][28] ),
    .A3(\core.cpuregs[27][28] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_05192_));
 sky130_fd_sc_hd__mux2_2 _11061_ (.A0(\core.cpuregs[30][28] ),
    .A1(\core.cpuregs[31][28] ),
    .S(_04437_),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_2 _11062_ (.A0(\core.cpuregs[28][28] ),
    .A1(\core.cpuregs[29][28] ),
    .S(_04600_),
    .X(_05194_));
 sky130_fd_sc_hd__a21o_2 _11063_ (.A1(_04512_),
    .A2(_05194_),
    .B1(_04526_),
    .X(_05195_));
 sky130_fd_sc_hd__a21o_2 _11064_ (.A1(_03326_),
    .A2(_05193_),
    .B1(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__o211a_2 _11065_ (.A1(_04519_),
    .A2(_05192_),
    .B1(_05196_),
    .C1(_03335_),
    .X(_05197_));
 sky130_fd_sc_hd__or3_2 _11066_ (.A(_04518_),
    .B(_05191_),
    .C(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__a32o_2 _11067_ (.A1(_04499_),
    .A2(_05185_),
    .A3(_05198_),
    .B1(_04541_),
    .B2(\core.reg_pc[28] ),
    .X(_05199_));
 sky130_fd_sc_hd__a22o_2 _11068_ (.A1(_02545_),
    .A2(_05172_),
    .B1(_05199_),
    .B2(_03261_),
    .X(_05200_));
 sky130_fd_sc_hd__a31o_2 _11069_ (.A1(_02042_),
    .A2(_05167_),
    .A3(_05168_),
    .B1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_2 _11070_ (.A0(_05201_),
    .A1(_02246_),
    .S(_04948_),
    .X(_05202_));
 sky130_fd_sc_hd__buf_1 _11071_ (.A(_05202_),
    .X(_00271_));
 sky130_fd_sc_hd__nor2_2 _11072_ (.A(_03348_),
    .B(_03349_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_2 _11073_ (.A(_03459_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__or2_2 _11074_ (.A(_03459_),
    .B(_05203_),
    .X(_05205_));
 sky130_fd_sc_hd__o21ai_2 _11075_ (.A1(_02814_),
    .A2(_04298_),
    .B1(_02099_),
    .Y(_05206_));
 sky130_fd_sc_hd__mux2_2 _11076_ (.A0(_02242_),
    .A1(_02246_),
    .S(_04613_),
    .X(_05207_));
 sky130_fd_sc_hd__a2bb2o_2 _11077_ (.A1_N(_05169_),
    .A2_N(_05206_),
    .B1(_05207_),
    .B2(_04575_),
    .X(_05208_));
 sky130_fd_sc_hd__mux4_2 _11078_ (.A0(\core.cpuregs[8][29] ),
    .A1(\core.cpuregs[9][29] ),
    .A2(\core.cpuregs[10][29] ),
    .A3(\core.cpuregs[11][29] ),
    .S0(_03296_),
    .S1(_03274_),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_2 _11079_ (.A0(\core.cpuregs[14][29] ),
    .A1(\core.cpuregs[15][29] ),
    .S(_03280_),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_2 _11080_ (.A0(\core.cpuregs[12][29] ),
    .A1(\core.cpuregs[13][29] ),
    .S(_03319_),
    .X(_05211_));
 sky130_fd_sc_hd__a21o_2 _11081_ (.A1(_03284_),
    .A2(_05211_),
    .B1(_03288_),
    .X(_05212_));
 sky130_fd_sc_hd__a21o_2 _11082_ (.A1(_04328_),
    .A2(_05210_),
    .B1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__o211a_2 _11083_ (.A1(_04325_),
    .A2(_05209_),
    .B1(_05213_),
    .C1(_04508_),
    .X(_05214_));
 sky130_fd_sc_hd__mux4_2 _11084_ (.A0(\core.cpuregs[4][29] ),
    .A1(\core.cpuregs[5][29] ),
    .A2(\core.cpuregs[6][29] ),
    .A3(\core.cpuregs[7][29] ),
    .S0(_04314_),
    .S1(_04583_),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_2 _11085_ (.A0(\core.cpuregs[2][29] ),
    .A1(\core.cpuregs[3][29] ),
    .S(_03304_),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_2 _11086_ (.A0(\core.cpuregs[0][29] ),
    .A1(\core.cpuregs[1][29] ),
    .S(_04524_),
    .X(_05217_));
 sky130_fd_sc_hd__a21o_2 _11087_ (.A1(_04523_),
    .A2(_05217_),
    .B1(_03267_),
    .X(_05218_));
 sky130_fd_sc_hd__a21o_2 _11088_ (.A1(_04521_),
    .A2(_05216_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__o211a_2 _11089_ (.A1(_03294_),
    .A2(_05215_),
    .B1(_05219_),
    .C1(_04529_),
    .X(_05220_));
 sky130_fd_sc_hd__or3_2 _11090_ (.A(_04500_),
    .B(_05214_),
    .C(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__mux4_2 _11091_ (.A0(\core.cpuregs[16][29] ),
    .A1(\core.cpuregs[17][29] ),
    .A2(\core.cpuregs[18][29] ),
    .A3(\core.cpuregs[19][29] ),
    .S0(_04431_),
    .S1(_03298_),
    .X(_05222_));
 sky130_fd_sc_hd__mux2_2 _11092_ (.A0(\core.cpuregs[22][29] ),
    .A1(\core.cpuregs[23][29] ),
    .S(_04592_),
    .X(_05223_));
 sky130_fd_sc_hd__mux2_2 _11093_ (.A0(\core.cpuregs[20][29] ),
    .A1(\core.cpuregs[21][29] ),
    .S(_03303_),
    .X(_05224_));
 sky130_fd_sc_hd__a21o_2 _11094_ (.A1(_04504_),
    .A2(_05224_),
    .B1(_03331_),
    .X(_05225_));
 sky130_fd_sc_hd__a21o_2 _11095_ (.A1(_04502_),
    .A2(_05223_),
    .B1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__o211a_2 _11096_ (.A1(_03315_),
    .A2(_05222_),
    .B1(_05226_),
    .C1(_03308_),
    .X(_05227_));
 sky130_fd_sc_hd__mux4_2 _11097_ (.A0(\core.cpuregs[24][29] ),
    .A1(\core.cpuregs[25][29] ),
    .A2(\core.cpuregs[26][29] ),
    .A3(\core.cpuregs[27][29] ),
    .S0(_04217_),
    .S1(_04433_),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_2 _11098_ (.A0(\core.cpuregs[30][29] ),
    .A1(\core.cpuregs[31][29] ),
    .S(_03329_),
    .X(_05229_));
 sky130_fd_sc_hd__mux2_2 _11099_ (.A0(\core.cpuregs[28][29] ),
    .A1(\core.cpuregs[29][29] ),
    .S(_04600_),
    .X(_05230_));
 sky130_fd_sc_hd__a21o_2 _11100_ (.A1(_04512_),
    .A2(_05230_),
    .B1(_04526_),
    .X(_05231_));
 sky130_fd_sc_hd__a21o_2 _11101_ (.A1(_03326_),
    .A2(_05229_),
    .B1(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__o211a_2 _11102_ (.A1(_04519_),
    .A2(_05228_),
    .B1(_05232_),
    .C1(_03335_),
    .X(_05233_));
 sky130_fd_sc_hd__or3_2 _11103_ (.A(_03312_),
    .B(_05227_),
    .C(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__a32o_2 _11104_ (.A1(_04499_),
    .A2(_05221_),
    .A3(_05234_),
    .B1(_04541_),
    .B2(\core.reg_pc[29] ),
    .X(_05235_));
 sky130_fd_sc_hd__a22o_2 _11105_ (.A1(_02545_),
    .A2(_05208_),
    .B1(_05235_),
    .B2(_03261_),
    .X(_05236_));
 sky130_fd_sc_hd__a31o_2 _11106_ (.A1(_02042_),
    .A2(_05204_),
    .A3(_05205_),
    .B1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_2 _11107_ (.A0(_05237_),
    .A1(_02414_),
    .S(_04948_),
    .X(_05238_));
 sky130_fd_sc_hd__buf_1 _11108_ (.A(_05238_),
    .X(_00272_));
 sky130_fd_sc_hd__a211o_2 _11109_ (.A1(_03347_),
    .A2(_03461_),
    .B1(_03348_),
    .C1(_03460_),
    .X(_05239_));
 sky130_fd_sc_hd__o21ba_2 _11110_ (.A1(_02422_),
    .A2(_04298_),
    .B1_N(_05169_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_2 _11111_ (.A0(_02237_),
    .A1(_02414_),
    .S(_04613_),
    .X(_05241_));
 sky130_fd_sc_hd__mux2_2 _11112_ (.A0(_05240_),
    .A1(_05241_),
    .S(_04575_),
    .X(_05242_));
 sky130_fd_sc_hd__a32o_2 _11113_ (.A1(_02041_),
    .A2(_03462_),
    .A3(_05239_),
    .B1(_05242_),
    .B2(_04244_),
    .X(_05243_));
 sky130_fd_sc_hd__mux4_2 _11114_ (.A0(\core.cpuregs[8][30] ),
    .A1(\core.cpuregs[9][30] ),
    .A2(\core.cpuregs[10][30] ),
    .A3(\core.cpuregs[11][30] ),
    .S0(_04218_),
    .S1(_04220_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_2 _11115_ (.A0(\core.cpuregs[14][30] ),
    .A1(\core.cpuregs[15][30] ),
    .S(_04385_),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_2 _11116_ (.A0(\core.cpuregs[12][30] ),
    .A1(\core.cpuregs[13][30] ),
    .S(_04326_),
    .X(_05246_));
 sky130_fd_sc_hd__a21o_2 _11117_ (.A1(_04404_),
    .A2(_05246_),
    .B1(_03332_),
    .X(_05247_));
 sky130_fd_sc_hd__a21o_2 _11118_ (.A1(_03327_),
    .A2(_05245_),
    .B1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__o211a_2 _11119_ (.A1(_03316_),
    .A2(_05244_),
    .B1(_05248_),
    .C1(_03336_),
    .X(_05249_));
 sky130_fd_sc_hd__mux4_2 _11120_ (.A0(\core.cpuregs[4][30] ),
    .A1(\core.cpuregs[5][30] ),
    .A2(\core.cpuregs[6][30] ),
    .A3(\core.cpuregs[7][30] ),
    .S0(_04255_),
    .S1(_04256_),
    .X(_05250_));
 sky130_fd_sc_hd__mux2_2 _11121_ (.A0(\core.cpuregs[2][30] ),
    .A1(\core.cpuregs[3][30] ),
    .S(_04446_),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_2 _11122_ (.A0(\core.cpuregs[0][30] ),
    .A1(\core.cpuregs[1][30] ),
    .S(_03272_),
    .X(_05252_));
 sky130_fd_sc_hd__a21o_2 _11123_ (.A1(_04469_),
    .A2(_05252_),
    .B1(_03268_),
    .X(_05253_));
 sky130_fd_sc_hd__a21o_2 _11124_ (.A1(_04467_),
    .A2(_05251_),
    .B1(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__o211a_2 _11125_ (.A1(_04260_),
    .A2(_05250_),
    .B1(_05254_),
    .C1(_04487_),
    .X(_05255_));
 sky130_fd_sc_hd__or3_2 _11126_ (.A(_03266_),
    .B(_05249_),
    .C(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__mux4_2 _11127_ (.A0(\core.cpuregs[28][30] ),
    .A1(\core.cpuregs[29][30] ),
    .A2(\core.cpuregs[30][30] ),
    .A3(\core.cpuregs[31][30] ),
    .S0(_04236_),
    .S1(_04237_),
    .X(_05257_));
 sky130_fd_sc_hd__mux4_2 _11128_ (.A0(\core.cpuregs[24][30] ),
    .A1(\core.cpuregs[25][30] ),
    .A2(\core.cpuregs[26][30] ),
    .A3(\core.cpuregs[27][30] ),
    .S0(_03297_),
    .S1(_03299_),
    .X(_05258_));
 sky130_fd_sc_hd__mux4_2 _11129_ (.A0(\core.cpuregs[20][30] ),
    .A1(\core.cpuregs[21][30] ),
    .A2(\core.cpuregs[22][30] ),
    .A3(\core.cpuregs[23][30] ),
    .S0(_04432_),
    .S1(_04434_),
    .X(_05259_));
 sky130_fd_sc_hd__mux4_2 _11130_ (.A0(\core.cpuregs[16][30] ),
    .A1(\core.cpuregs[17][30] ),
    .A2(\core.cpuregs[18][30] ),
    .A3(\core.cpuregs[19][30] ),
    .S0(_04399_),
    .S1(_04400_),
    .X(_05260_));
 sky130_fd_sc_hd__mux4_2 _11131_ (.A0(_05257_),
    .A1(_05258_),
    .A2(_05259_),
    .A3(_05260_),
    .S0(_04266_),
    .S1(_04409_),
    .X(_05261_));
 sky130_fd_sc_hd__o21a_2 _11132_ (.A1(_03313_),
    .A2(_05261_),
    .B1(_04293_),
    .X(_05262_));
 sky130_fd_sc_hd__a221o_2 _11133_ (.A1(\core.reg_pc[30] ),
    .A2(_04253_),
    .B1(_05256_),
    .B2(_05262_),
    .C1(_04490_),
    .X(_05263_));
 sky130_fd_sc_hd__o21a_2 _11134_ (.A1(_03262_),
    .A2(_05243_),
    .B1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__mux2_2 _11135_ (.A0(_05264_),
    .A1(_02242_),
    .S(_03473_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_1 _11136_ (.A(_05265_),
    .X(_00273_));
 sky130_fd_sc_hd__or2_2 _11137_ (.A(\core.mem_do_wdata ),
    .B(_02027_),
    .X(_05266_));
 sky130_fd_sc_hd__or4b_2 _11138_ (.A(\core.mem_do_rinst ),
    .B(\core.mem_do_rdata ),
    .C(\core.mem_state[1] ),
    .D_N(\core.mem_state[0] ),
    .X(_05267_));
 sky130_fd_sc_hd__or2_2 _11139_ (.A(_02048_),
    .B(trap),
    .X(_05268_));
 sky130_fd_sc_hd__buf_1 _11140_ (.A(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__a21oi_2 _11141_ (.A1(_05266_),
    .A2(_05267_),
    .B1(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_2 _11142_ (.A(\core.mem_state[1] ),
    .B(\core.mem_state[0] ),
    .Y(_05271_));
 sky130_fd_sc_hd__or4b_2 _11143_ (.A(_03176_),
    .B(_05268_),
    .C(_03209_),
    .D_N(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__o41a_2 _11144_ (.A1(\core.mem_do_rdata ),
    .A2(_03206_),
    .A3(_05268_),
    .A4(_05266_),
    .B1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__nand2_2 _11145_ (.A(_02024_),
    .B(trap),
    .Y(_05274_));
 sky130_fd_sc_hd__o311a_2 _11146_ (.A1(\core.mem_do_rinst ),
    .A2(_05271_),
    .A3(_05269_),
    .B1(_05273_),
    .C1(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__mux2_2 _11147_ (.A0(\core.mem_state[0] ),
    .A1(_05270_),
    .S(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__buf_1 _11148_ (.A(_05276_),
    .X(_00274_));
 sky130_fd_sc_hd__a21oi_2 _11149_ (.A1(_03211_),
    .A2(_05267_),
    .B1(_05269_),
    .Y(_05277_));
 sky130_fd_sc_hd__mux2_2 _11150_ (.A0(\core.mem_state[1] ),
    .A1(_05277_),
    .S(_05275_),
    .X(_05278_));
 sky130_fd_sc_hd__buf_1 _11151_ (.A(_05278_),
    .X(_00275_));
 sky130_fd_sc_hd__and2b_2 _11152_ (.A_N(\core.latched_branch ),
    .B(\core.latched_store ),
    .X(_05279_));
 sky130_fd_sc_hd__buf_1 _11153_ (.A(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__buf_1 _11154_ (.A(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__mux2_2 _11155_ (.A0(\core.reg_out[0] ),
    .A1(\core.alu_out_q[0] ),
    .S(_03862_),
    .X(_05282_));
 sky130_fd_sc_hd__and2_2 _11156_ (.A(_05281_),
    .B(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__buf_1 _11157_ (.A(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__nand3b_2 _11158_ (.A_N(\core.latched_rd[3] ),
    .B(\core.latched_rd[2] ),
    .C(\core.latched_rd[4] ),
    .Y(_05285_));
 sky130_fd_sc_hd__o2111ai_2 _11159_ (.A1(\core.latched_store ),
    .A2(\core.latched_branch ),
    .B1(\core.latched_rd[1] ),
    .C1(\core.latched_rd[0] ),
    .D1(_02111_),
    .Y(_05286_));
 sky130_fd_sc_hd__nor2_2 _11160_ (.A(_05285_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__buf_1 _11161_ (.A(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_2 _11162_ (.A0(\core.cpuregs[23][0] ),
    .A1(_05284_),
    .S(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__buf_1 _11163_ (.A(_05289_),
    .X(_00276_));
 sky130_fd_sc_hd__buf_1 _11164_ (.A(_05280_),
    .X(_05290_));
 sky130_fd_sc_hd__mux2_2 _11165_ (.A0(\core.reg_pc[1] ),
    .A1(_03657_),
    .S(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__buf_1 _11166_ (.A(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__mux2_2 _11167_ (.A0(\core.cpuregs[23][1] ),
    .A1(_05292_),
    .S(_05288_),
    .X(_05293_));
 sky130_fd_sc_hd__buf_1 _11168_ (.A(_05293_),
    .X(_00277_));
 sky130_fd_sc_hd__inv_2 _11169_ (.A(_02493_),
    .Y(_05294_));
 sky130_fd_sc_hd__buf_1 _11170_ (.A(_05280_),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_2 _11171_ (.A0(_05294_),
    .A1(_03668_),
    .S(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__buf_1 _11172_ (.A(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__mux2_2 _11173_ (.A0(\core.cpuregs[23][2] ),
    .A1(_05297_),
    .S(_05288_),
    .X(_05298_));
 sky130_fd_sc_hd__buf_1 _11174_ (.A(_05298_),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_2 _11175_ (.A(\core.reg_pc[3] ),
    .B(_02493_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2b_2 _11176_ (.A_N(\core.latched_branch ),
    .B(\core.latched_store ),
    .Y(_05300_));
 sky130_fd_sc_hd__buf_1 _11177_ (.A(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__o21a_2 _11178_ (.A1(\core.reg_pc[3] ),
    .A2(_02493_),
    .B1(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__a22o_2 _11179_ (.A1(_03682_),
    .A2(_05281_),
    .B1(_05299_),
    .B2(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__buf_1 _11180_ (.A(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_2 _11181_ (.A0(\core.cpuregs[23][3] ),
    .A1(_05304_),
    .S(_05288_),
    .X(_05305_));
 sky130_fd_sc_hd__buf_1 _11182_ (.A(_05305_),
    .X(_00279_));
 sky130_fd_sc_hd__a21o_2 _11183_ (.A1(\core.reg_pc[3] ),
    .A2(_02493_),
    .B1(\core.reg_pc[4] ),
    .X(_05306_));
 sky130_fd_sc_hd__and3_2 _11184_ (.A(\core.reg_pc[4] ),
    .B(\core.reg_pc[3] ),
    .C(_02493_),
    .X(_05307_));
 sky130_fd_sc_hd__nor2_2 _11185_ (.A(_05295_),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__a22o_2 _11186_ (.A1(_03700_),
    .A2(_05281_),
    .B1(_05306_),
    .B2(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__buf_1 _11187_ (.A(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__mux2_2 _11188_ (.A0(\core.cpuregs[23][4] ),
    .A1(_05310_),
    .S(_05288_),
    .X(_05311_));
 sky130_fd_sc_hd__buf_1 _11189_ (.A(_05311_),
    .X(_00280_));
 sky130_fd_sc_hd__o21ai_2 _11190_ (.A1(\core.reg_pc[5] ),
    .A2(_05307_),
    .B1(_05301_),
    .Y(_05312_));
 sky130_fd_sc_hd__and4_2 _11191_ (.A(\core.reg_pc[5] ),
    .B(\core.reg_pc[4] ),
    .C(\core.reg_pc[3] ),
    .D(\core.reg_pc[2] ),
    .X(_05313_));
 sky130_fd_sc_hd__a2bb2o_2 _11192_ (.A1_N(_05312_),
    .A2_N(_05313_),
    .B1(_05290_),
    .B2(_03716_),
    .X(_05314_));
 sky130_fd_sc_hd__buf_1 _11193_ (.A(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__mux2_2 _11194_ (.A0(\core.cpuregs[23][5] ),
    .A1(_05315_),
    .S(_05288_),
    .X(_05316_));
 sky130_fd_sc_hd__buf_1 _11195_ (.A(_05316_),
    .X(_00281_));
 sky130_fd_sc_hd__or2_2 _11196_ (.A(\core.reg_pc[6] ),
    .B(_05313_),
    .X(_05317_));
 sky130_fd_sc_hd__a21oi_2 _11197_ (.A1(\core.reg_pc[6] ),
    .A2(_05313_),
    .B1(_05295_),
    .Y(_05318_));
 sky130_fd_sc_hd__a22o_2 _11198_ (.A1(_03730_),
    .A2(_05281_),
    .B1(_05317_),
    .B2(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__buf_1 _11199_ (.A(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_2 _11200_ (.A0(\core.cpuregs[23][6] ),
    .A1(_05320_),
    .S(_05288_),
    .X(_05321_));
 sky130_fd_sc_hd__buf_1 _11201_ (.A(_05321_),
    .X(_00282_));
 sky130_fd_sc_hd__a21oi_2 _11202_ (.A1(\core.reg_pc[6] ),
    .A2(_05313_),
    .B1(\core.reg_pc[7] ),
    .Y(_05322_));
 sky130_fd_sc_hd__and3_2 _11203_ (.A(\core.reg_pc[7] ),
    .B(\core.reg_pc[6] ),
    .C(_05313_),
    .X(_05323_));
 sky130_fd_sc_hd__nor2_2 _11204_ (.A(_05322_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__mux2_2 _11205_ (.A0(_03740_),
    .A1(_05324_),
    .S(_05301_),
    .X(_05325_));
 sky130_fd_sc_hd__buf_1 _11206_ (.A(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_2 _11207_ (.A0(\core.cpuregs[23][7] ),
    .A1(_05326_),
    .S(_05288_),
    .X(_05327_));
 sky130_fd_sc_hd__buf_1 _11208_ (.A(_05327_),
    .X(_00283_));
 sky130_fd_sc_hd__or2_2 _11209_ (.A(\core.reg_pc[8] ),
    .B(_05323_),
    .X(_05328_));
 sky130_fd_sc_hd__and4_2 _11210_ (.A(\core.reg_pc[8] ),
    .B(\core.reg_pc[7] ),
    .C(\core.reg_pc[6] ),
    .D(_05313_),
    .X(_05329_));
 sky130_fd_sc_hd__nor2_2 _11211_ (.A(_05295_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__a22o_2 _11212_ (.A1(_03751_),
    .A2(_05281_),
    .B1(_05328_),
    .B2(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__buf_1 _11213_ (.A(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_2 _11214_ (.A0(\core.cpuregs[23][8] ),
    .A1(_05332_),
    .S(_05288_),
    .X(_05333_));
 sky130_fd_sc_hd__buf_1 _11215_ (.A(_05333_),
    .X(_00284_));
 sky130_fd_sc_hd__nand2_2 _11216_ (.A(\core.reg_pc[9] ),
    .B(_05329_),
    .Y(_05334_));
 sky130_fd_sc_hd__o21a_2 _11217_ (.A1(\core.reg_pc[9] ),
    .A2(_05329_),
    .B1(_05301_),
    .X(_05335_));
 sky130_fd_sc_hd__a22o_2 _11218_ (.A1(_03770_),
    .A2(_05281_),
    .B1(_05334_),
    .B2(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__buf_1 _11219_ (.A(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_2 _11220_ (.A0(\core.cpuregs[23][9] ),
    .A1(_05337_),
    .S(_05288_),
    .X(_05338_));
 sky130_fd_sc_hd__buf_1 _11221_ (.A(_05338_),
    .X(_00285_));
 sky130_fd_sc_hd__a21o_2 _11222_ (.A1(\core.reg_pc[9] ),
    .A2(_05329_),
    .B1(\core.reg_pc[10] ),
    .X(_05339_));
 sky130_fd_sc_hd__and3_2 _11223_ (.A(\core.reg_pc[10] ),
    .B(\core.reg_pc[9] ),
    .C(_05329_),
    .X(_05340_));
 sky130_fd_sc_hd__nor2_2 _11224_ (.A(_05295_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__a22o_2 _11225_ (.A1(_03781_),
    .A2(_05281_),
    .B1(_05339_),
    .B2(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__buf_1 _11226_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__buf_1 _11227_ (.A(_05287_),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_2 _11228_ (.A0(\core.cpuregs[23][10] ),
    .A1(_05343_),
    .S(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__buf_1 _11229_ (.A(_05345_),
    .X(_00286_));
 sky130_fd_sc_hd__or2_2 _11230_ (.A(\core.reg_pc[11] ),
    .B(_05340_),
    .X(_05346_));
 sky130_fd_sc_hd__a21oi_2 _11231_ (.A1(\core.reg_pc[11] ),
    .A2(_05340_),
    .B1(_05295_),
    .Y(_05347_));
 sky130_fd_sc_hd__a22o_2 _11232_ (.A1(_03794_),
    .A2(_05281_),
    .B1(_05346_),
    .B2(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__buf_1 _11233_ (.A(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_2 _11234_ (.A0(\core.cpuregs[23][11] ),
    .A1(_05349_),
    .S(_05344_),
    .X(_05350_));
 sky130_fd_sc_hd__buf_1 _11235_ (.A(_05350_),
    .X(_00287_));
 sky130_fd_sc_hd__a21o_2 _11236_ (.A1(\core.reg_pc[11] ),
    .A2(_05340_),
    .B1(\core.reg_pc[12] ),
    .X(_05351_));
 sky130_fd_sc_hd__and3_2 _11237_ (.A(\core.reg_pc[12] ),
    .B(\core.reg_pc[11] ),
    .C(_05340_),
    .X(_05352_));
 sky130_fd_sc_hd__nor2_2 _11238_ (.A(_05295_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__a22o_2 _11239_ (.A1(_03806_),
    .A2(_05281_),
    .B1(_05351_),
    .B2(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__buf_1 _11240_ (.A(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_2 _11241_ (.A0(\core.cpuregs[23][12] ),
    .A1(_05355_),
    .S(_05344_),
    .X(_05356_));
 sky130_fd_sc_hd__buf_1 _11242_ (.A(_05356_),
    .X(_00288_));
 sky130_fd_sc_hd__or2_2 _11243_ (.A(\core.reg_pc[13] ),
    .B(_05352_),
    .X(_05357_));
 sky130_fd_sc_hd__a21oi_2 _11244_ (.A1(\core.reg_pc[13] ),
    .A2(_05352_),
    .B1(_05295_),
    .Y(_05358_));
 sky130_fd_sc_hd__a22o_2 _11245_ (.A1(_03825_),
    .A2(_05281_),
    .B1(_05357_),
    .B2(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__buf_1 _11246_ (.A(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_2 _11247_ (.A0(\core.cpuregs[23][13] ),
    .A1(_05360_),
    .S(_05344_),
    .X(_05361_));
 sky130_fd_sc_hd__buf_1 _11248_ (.A(_05361_),
    .X(_00289_));
 sky130_fd_sc_hd__buf_1 _11249_ (.A(_05280_),
    .X(_05362_));
 sky130_fd_sc_hd__a21o_2 _11250_ (.A1(\core.reg_pc[13] ),
    .A2(_05352_),
    .B1(\core.reg_pc[14] ),
    .X(_05363_));
 sky130_fd_sc_hd__and3_2 _11251_ (.A(\core.reg_pc[14] ),
    .B(\core.reg_pc[13] ),
    .C(_05352_),
    .X(_05364_));
 sky130_fd_sc_hd__nor2_2 _11252_ (.A(_05280_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__a22o_2 _11253_ (.A1(_03836_),
    .A2(_05362_),
    .B1(_05363_),
    .B2(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__buf_1 _11254_ (.A(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_2 _11255_ (.A0(\core.cpuregs[23][14] ),
    .A1(_05367_),
    .S(_05344_),
    .X(_05368_));
 sky130_fd_sc_hd__buf_1 _11256_ (.A(_05368_),
    .X(_00290_));
 sky130_fd_sc_hd__o21ai_2 _11257_ (.A1(\core.reg_pc[15] ),
    .A2(_05364_),
    .B1(_05301_),
    .Y(_05369_));
 sky130_fd_sc_hd__and2_2 _11258_ (.A(\core.reg_pc[15] ),
    .B(_05364_),
    .X(_05370_));
 sky130_fd_sc_hd__a2bb2o_2 _11259_ (.A1_N(_05369_),
    .A2_N(_05370_),
    .B1(_05290_),
    .B2(_03847_),
    .X(_05371_));
 sky130_fd_sc_hd__buf_1 _11260_ (.A(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__mux2_2 _11261_ (.A0(\core.cpuregs[23][15] ),
    .A1(_05372_),
    .S(_05344_),
    .X(_05373_));
 sky130_fd_sc_hd__buf_1 _11262_ (.A(_05373_),
    .X(_00291_));
 sky130_fd_sc_hd__or2_2 _11263_ (.A(\core.reg_pc[16] ),
    .B(_05370_),
    .X(_05374_));
 sky130_fd_sc_hd__a21oi_2 _11264_ (.A1(\core.reg_pc[16] ),
    .A2(_05370_),
    .B1(_05295_),
    .Y(_05375_));
 sky130_fd_sc_hd__a22o_2 _11265_ (.A1(_03863_),
    .A2(_05362_),
    .B1(_05374_),
    .B2(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__buf_1 _11266_ (.A(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__mux2_2 _11267_ (.A0(\core.cpuregs[23][16] ),
    .A1(_05377_),
    .S(_05344_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_1 _11268_ (.A(_05378_),
    .X(_00292_));
 sky130_fd_sc_hd__a31o_2 _11269_ (.A1(\core.reg_pc[16] ),
    .A2(\core.reg_pc[15] ),
    .A3(_05364_),
    .B1(\core.reg_pc[17] ),
    .X(_05379_));
 sky130_fd_sc_hd__and3_2 _11270_ (.A(\core.reg_pc[17] ),
    .B(\core.reg_pc[16] ),
    .C(_05370_),
    .X(_05380_));
 sky130_fd_sc_hd__nor2_2 _11271_ (.A(_05280_),
    .B(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__a22o_2 _11272_ (.A1(_03881_),
    .A2(_05362_),
    .B1(_05379_),
    .B2(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__buf_1 _11273_ (.A(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__mux2_2 _11274_ (.A0(\core.cpuregs[23][17] ),
    .A1(_05383_),
    .S(_05344_),
    .X(_05384_));
 sky130_fd_sc_hd__buf_1 _11275_ (.A(_05384_),
    .X(_00293_));
 sky130_fd_sc_hd__o21ai_2 _11276_ (.A1(\core.reg_pc[18] ),
    .A2(_05380_),
    .B1(_05301_),
    .Y(_05385_));
 sky130_fd_sc_hd__and2_2 _11277_ (.A(\core.reg_pc[18] ),
    .B(_05380_),
    .X(_05386_));
 sky130_fd_sc_hd__a2bb2o_2 _11278_ (.A1_N(_05385_),
    .A2_N(_05386_),
    .B1(_05290_),
    .B2(_03892_),
    .X(_05387_));
 sky130_fd_sc_hd__buf_1 _11279_ (.A(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__mux2_2 _11280_ (.A0(\core.cpuregs[23][18] ),
    .A1(_05388_),
    .S(_05344_),
    .X(_05389_));
 sky130_fd_sc_hd__buf_1 _11281_ (.A(_05389_),
    .X(_00294_));
 sky130_fd_sc_hd__nand2_2 _11282_ (.A(\core.reg_pc[19] ),
    .B(_05386_),
    .Y(_05390_));
 sky130_fd_sc_hd__o21a_2 _11283_ (.A1(\core.reg_pc[19] ),
    .A2(_05386_),
    .B1(_05300_),
    .X(_05391_));
 sky130_fd_sc_hd__a22o_2 _11284_ (.A1(_03902_),
    .A2(_05362_),
    .B1(_05390_),
    .B2(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__buf_1 _11285_ (.A(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__mux2_2 _11286_ (.A0(\core.cpuregs[23][19] ),
    .A1(_05393_),
    .S(_05344_),
    .X(_05394_));
 sky130_fd_sc_hd__buf_1 _11287_ (.A(_05394_),
    .X(_00295_));
 sky130_fd_sc_hd__a31o_2 _11288_ (.A1(\core.reg_pc[19] ),
    .A2(\core.reg_pc[18] ),
    .A3(_05380_),
    .B1(\core.reg_pc[20] ),
    .X(_05395_));
 sky130_fd_sc_hd__and3_2 _11289_ (.A(\core.reg_pc[20] ),
    .B(\core.reg_pc[19] ),
    .C(_05386_),
    .X(_05396_));
 sky130_fd_sc_hd__nor2_2 _11290_ (.A(_05280_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a22o_2 _11291_ (.A1(_03916_),
    .A2(_05362_),
    .B1(_05395_),
    .B2(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__buf_1 _11292_ (.A(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__buf_1 _11293_ (.A(_05287_),
    .X(_05400_));
 sky130_fd_sc_hd__mux2_2 _11294_ (.A0(\core.cpuregs[23][20] ),
    .A1(_05399_),
    .S(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__buf_1 _11295_ (.A(_05401_),
    .X(_00296_));
 sky130_fd_sc_hd__o21ai_2 _11296_ (.A1(\core.reg_pc[21] ),
    .A2(_05396_),
    .B1(_05301_),
    .Y(_05402_));
 sky130_fd_sc_hd__and2_2 _11297_ (.A(\core.reg_pc[21] ),
    .B(_05396_),
    .X(_05403_));
 sky130_fd_sc_hd__a2bb2o_2 _11298_ (.A1_N(_05402_),
    .A2_N(_05403_),
    .B1(_05290_),
    .B2(_03928_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_1 _11299_ (.A(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_2 _11300_ (.A0(\core.cpuregs[23][21] ),
    .A1(_05405_),
    .S(_05400_),
    .X(_05406_));
 sky130_fd_sc_hd__buf_1 _11301_ (.A(_05406_),
    .X(_00297_));
 sky130_fd_sc_hd__nand2_2 _11302_ (.A(\core.reg_pc[22] ),
    .B(_05403_),
    .Y(_05407_));
 sky130_fd_sc_hd__o21a_2 _11303_ (.A1(\core.reg_pc[22] ),
    .A2(_05403_),
    .B1(_05300_),
    .X(_05408_));
 sky130_fd_sc_hd__a22o_2 _11304_ (.A1(_03945_),
    .A2(_05362_),
    .B1(_05407_),
    .B2(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__buf_1 _11305_ (.A(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__mux2_2 _11306_ (.A0(\core.cpuregs[23][22] ),
    .A1(_05410_),
    .S(_05400_),
    .X(_05411_));
 sky130_fd_sc_hd__buf_1 _11307_ (.A(_05411_),
    .X(_00298_));
 sky130_fd_sc_hd__a31o_2 _11308_ (.A1(\core.reg_pc[22] ),
    .A2(\core.reg_pc[21] ),
    .A3(_05396_),
    .B1(\core.reg_pc[23] ),
    .X(_05412_));
 sky130_fd_sc_hd__and3_2 _11309_ (.A(\core.reg_pc[23] ),
    .B(\core.reg_pc[22] ),
    .C(_05403_),
    .X(_05413_));
 sky130_fd_sc_hd__nor2_2 _11310_ (.A(_05280_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__a22o_2 _11311_ (.A1(_03956_),
    .A2(_05362_),
    .B1(_05412_),
    .B2(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__buf_1 _11312_ (.A(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__mux2_2 _11313_ (.A0(\core.cpuregs[23][23] ),
    .A1(_05416_),
    .S(_05400_),
    .X(_05417_));
 sky130_fd_sc_hd__buf_1 _11314_ (.A(_05417_),
    .X(_00299_));
 sky130_fd_sc_hd__o21ai_2 _11315_ (.A1(\core.reg_pc[24] ),
    .A2(_05413_),
    .B1(_05301_),
    .Y(_05418_));
 sky130_fd_sc_hd__and2_2 _11316_ (.A(\core.reg_pc[24] ),
    .B(_05413_),
    .X(_05419_));
 sky130_fd_sc_hd__a2bb2o_2 _11317_ (.A1_N(_05418_),
    .A2_N(_05419_),
    .B1(_05290_),
    .B2(_03971_),
    .X(_05420_));
 sky130_fd_sc_hd__buf_1 _11318_ (.A(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_2 _11319_ (.A0(\core.cpuregs[23][24] ),
    .A1(_05421_),
    .S(_05400_),
    .X(_05422_));
 sky130_fd_sc_hd__buf_1 _11320_ (.A(_05422_),
    .X(_00300_));
 sky130_fd_sc_hd__nand2_2 _11321_ (.A(\core.reg_pc[25] ),
    .B(_05419_),
    .Y(_05423_));
 sky130_fd_sc_hd__o21a_2 _11322_ (.A1(\core.reg_pc[25] ),
    .A2(_05419_),
    .B1(_05300_),
    .X(_05424_));
 sky130_fd_sc_hd__a22o_2 _11323_ (.A1(_03988_),
    .A2(_05362_),
    .B1(_05423_),
    .B2(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__buf_1 _11324_ (.A(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_2 _11325_ (.A0(\core.cpuregs[23][25] ),
    .A1(_05426_),
    .S(_05400_),
    .X(_05427_));
 sky130_fd_sc_hd__buf_1 _11326_ (.A(_05427_),
    .X(_00301_));
 sky130_fd_sc_hd__a31o_2 _11327_ (.A1(\core.reg_pc[25] ),
    .A2(\core.reg_pc[24] ),
    .A3(_05413_),
    .B1(\core.reg_pc[26] ),
    .X(_05428_));
 sky130_fd_sc_hd__and3_2 _11328_ (.A(\core.reg_pc[26] ),
    .B(\core.reg_pc[25] ),
    .C(_05419_),
    .X(_05429_));
 sky130_fd_sc_hd__nor2_2 _11329_ (.A(_05280_),
    .B(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__a22o_2 _11330_ (.A1(_03997_),
    .A2(_05362_),
    .B1(_05428_),
    .B2(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__buf_1 _11331_ (.A(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_2 _11332_ (.A0(\core.cpuregs[23][26] ),
    .A1(_05432_),
    .S(_05400_),
    .X(_05433_));
 sky130_fd_sc_hd__buf_1 _11333_ (.A(_05433_),
    .X(_00302_));
 sky130_fd_sc_hd__o21ai_2 _11334_ (.A1(\core.reg_pc[27] ),
    .A2(_05429_),
    .B1(_05301_),
    .Y(_05434_));
 sky130_fd_sc_hd__and2_2 _11335_ (.A(\core.reg_pc[27] ),
    .B(_05429_),
    .X(_05435_));
 sky130_fd_sc_hd__a2bb2o_2 _11336_ (.A1_N(_05434_),
    .A2_N(_05435_),
    .B1(_05290_),
    .B2(_04010_),
    .X(_05436_));
 sky130_fd_sc_hd__buf_1 _11337_ (.A(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_2 _11338_ (.A0(\core.cpuregs[23][27] ),
    .A1(_05437_),
    .S(_05400_),
    .X(_05438_));
 sky130_fd_sc_hd__buf_1 _11339_ (.A(_05438_),
    .X(_00303_));
 sky130_fd_sc_hd__or2_2 _11340_ (.A(\core.reg_pc[28] ),
    .B(_05435_),
    .X(_05439_));
 sky130_fd_sc_hd__a21oi_2 _11341_ (.A1(\core.reg_pc[28] ),
    .A2(_05435_),
    .B1(_05295_),
    .Y(_05440_));
 sky130_fd_sc_hd__a22o_2 _11342_ (.A1(_04019_),
    .A2(_05362_),
    .B1(_05439_),
    .B2(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__buf_1 _11343_ (.A(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__mux2_2 _11344_ (.A0(\core.cpuregs[23][28] ),
    .A1(_05442_),
    .S(_05400_),
    .X(_05443_));
 sky130_fd_sc_hd__buf_1 _11345_ (.A(_05443_),
    .X(_00304_));
 sky130_fd_sc_hd__a31o_2 _11346_ (.A1(\core.reg_pc[28] ),
    .A2(\core.reg_pc[27] ),
    .A3(_05429_),
    .B1(\core.reg_pc[29] ),
    .X(_05444_));
 sky130_fd_sc_hd__and3_2 _11347_ (.A(\core.reg_pc[29] ),
    .B(\core.reg_pc[28] ),
    .C(_05435_),
    .X(_05445_));
 sky130_fd_sc_hd__nor2_2 _11348_ (.A(_05280_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__a22o_2 _11349_ (.A1(_04031_),
    .A2(_05290_),
    .B1(_05444_),
    .B2(_05446_),
    .X(_05447_));
 sky130_fd_sc_hd__buf_1 _11350_ (.A(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__mux2_2 _11351_ (.A0(\core.cpuregs[23][29] ),
    .A1(_05448_),
    .S(_05400_),
    .X(_05449_));
 sky130_fd_sc_hd__buf_1 _11352_ (.A(_05449_),
    .X(_00305_));
 sky130_fd_sc_hd__o21ai_2 _11353_ (.A1(\core.reg_pc[30] ),
    .A2(_05445_),
    .B1(_05301_),
    .Y(_05450_));
 sky130_fd_sc_hd__and2_2 _11354_ (.A(\core.reg_pc[30] ),
    .B(_05445_),
    .X(_05451_));
 sky130_fd_sc_hd__a2bb2o_2 _11355_ (.A1_N(_05450_),
    .A2_N(_05451_),
    .B1(_05290_),
    .B2(_04041_),
    .X(_05452_));
 sky130_fd_sc_hd__buf_1 _11356_ (.A(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__mux2_2 _11357_ (.A0(\core.cpuregs[23][30] ),
    .A1(_05453_),
    .S(_05287_),
    .X(_05454_));
 sky130_fd_sc_hd__buf_1 _11358_ (.A(_05454_),
    .X(_00306_));
 sky130_fd_sc_hd__nand2_2 _11359_ (.A(\core.reg_pc[31] ),
    .B(_05451_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21a_2 _11360_ (.A1(\core.reg_pc[31] ),
    .A2(_05451_),
    .B1(_05300_),
    .X(_05456_));
 sky130_fd_sc_hd__a22o_2 _11361_ (.A1(_04053_),
    .A2(_05290_),
    .B1(_05455_),
    .B2(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__buf_1 _11362_ (.A(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__mux2_2 _11363_ (.A0(\core.cpuregs[23][31] ),
    .A1(_05458_),
    .S(_05287_),
    .X(_05459_));
 sky130_fd_sc_hd__buf_1 _11364_ (.A(_05459_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_1 _11365_ (.A(_05283_),
    .X(_05460_));
 sky130_fd_sc_hd__nand3_2 _11366_ (.A(\core.latched_rd[4] ),
    .B(\core.latched_rd[3] ),
    .C(\core.latched_rd[2] ),
    .Y(_05461_));
 sky130_fd_sc_hd__o21ai_2 _11367_ (.A1(\core.latched_store ),
    .A2(\core.latched_branch ),
    .B1(_02111_),
    .Y(_05462_));
 sky130_fd_sc_hd__or3b_2 _11368_ (.A(\core.latched_rd[0] ),
    .B(_05462_),
    .C_N(\core.latched_rd[1] ),
    .X(_05463_));
 sky130_fd_sc_hd__buf_1 _11369_ (.A(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__or2_2 _11370_ (.A(_05461_),
    .B(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__buf_1 _11371_ (.A(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_2 _11372_ (.A0(_05460_),
    .A1(\core.cpuregs[30][0] ),
    .S(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__buf_1 _11373_ (.A(_05467_),
    .X(_00308_));
 sky130_fd_sc_hd__buf_1 _11374_ (.A(_05291_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_2 _11375_ (.A0(_05468_),
    .A1(\core.cpuregs[30][1] ),
    .S(_05466_),
    .X(_05469_));
 sky130_fd_sc_hd__buf_1 _11376_ (.A(_05469_),
    .X(_00309_));
 sky130_fd_sc_hd__buf_1 _11377_ (.A(_05296_),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_2 _11378_ (.A0(_05470_),
    .A1(\core.cpuregs[30][2] ),
    .S(_05466_),
    .X(_05471_));
 sky130_fd_sc_hd__buf_1 _11379_ (.A(_05471_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_1 _11380_ (.A(_05303_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_2 _11381_ (.A0(_05472_),
    .A1(\core.cpuregs[30][3] ),
    .S(_05466_),
    .X(_05473_));
 sky130_fd_sc_hd__buf_1 _11382_ (.A(_05473_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_1 _11383_ (.A(_05309_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_2 _11384_ (.A0(_05474_),
    .A1(\core.cpuregs[30][4] ),
    .S(_05466_),
    .X(_05475_));
 sky130_fd_sc_hd__buf_1 _11385_ (.A(_05475_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_1 _11386_ (.A(_05314_),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_2 _11387_ (.A0(_05476_),
    .A1(\core.cpuregs[30][5] ),
    .S(_05466_),
    .X(_05477_));
 sky130_fd_sc_hd__buf_1 _11388_ (.A(_05477_),
    .X(_00313_));
 sky130_fd_sc_hd__buf_1 _11389_ (.A(_05319_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_2 _11390_ (.A0(_05478_),
    .A1(\core.cpuregs[30][6] ),
    .S(_05466_),
    .X(_05479_));
 sky130_fd_sc_hd__buf_1 _11391_ (.A(_05479_),
    .X(_00314_));
 sky130_fd_sc_hd__buf_1 _11392_ (.A(_05325_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_2 _11393_ (.A0(_05480_),
    .A1(\core.cpuregs[30][7] ),
    .S(_05466_),
    .X(_05481_));
 sky130_fd_sc_hd__buf_1 _11394_ (.A(_05481_),
    .X(_00315_));
 sky130_fd_sc_hd__buf_1 _11395_ (.A(_05331_),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_2 _11396_ (.A0(_05482_),
    .A1(\core.cpuregs[30][8] ),
    .S(_05466_),
    .X(_05483_));
 sky130_fd_sc_hd__buf_1 _11397_ (.A(_05483_),
    .X(_00316_));
 sky130_fd_sc_hd__buf_1 _11398_ (.A(_05336_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_2 _11399_ (.A0(_05484_),
    .A1(\core.cpuregs[30][9] ),
    .S(_05466_),
    .X(_05485_));
 sky130_fd_sc_hd__buf_1 _11400_ (.A(_05485_),
    .X(_00317_));
 sky130_fd_sc_hd__buf_1 _11401_ (.A(_05342_),
    .X(_05486_));
 sky130_fd_sc_hd__buf_1 _11402_ (.A(_05465_),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_2 _11403_ (.A0(_05486_),
    .A1(\core.cpuregs[30][10] ),
    .S(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__buf_1 _11404_ (.A(_05488_),
    .X(_00318_));
 sky130_fd_sc_hd__buf_1 _11405_ (.A(_05348_),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_2 _11406_ (.A0(_05489_),
    .A1(\core.cpuregs[30][11] ),
    .S(_05487_),
    .X(_05490_));
 sky130_fd_sc_hd__buf_1 _11407_ (.A(_05490_),
    .X(_00319_));
 sky130_fd_sc_hd__buf_1 _11408_ (.A(_05354_),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_2 _11409_ (.A0(_05491_),
    .A1(\core.cpuregs[30][12] ),
    .S(_05487_),
    .X(_05492_));
 sky130_fd_sc_hd__buf_1 _11410_ (.A(_05492_),
    .X(_00320_));
 sky130_fd_sc_hd__buf_1 _11411_ (.A(_05359_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_2 _11412_ (.A0(_05493_),
    .A1(\core.cpuregs[30][13] ),
    .S(_05487_),
    .X(_05494_));
 sky130_fd_sc_hd__buf_1 _11413_ (.A(_05494_),
    .X(_00321_));
 sky130_fd_sc_hd__buf_1 _11414_ (.A(_05366_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_2 _11415_ (.A0(_05495_),
    .A1(\core.cpuregs[30][14] ),
    .S(_05487_),
    .X(_05496_));
 sky130_fd_sc_hd__buf_1 _11416_ (.A(_05496_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_1 _11417_ (.A(_05371_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_2 _11418_ (.A0(_05497_),
    .A1(\core.cpuregs[30][15] ),
    .S(_05487_),
    .X(_05498_));
 sky130_fd_sc_hd__buf_1 _11419_ (.A(_05498_),
    .X(_00323_));
 sky130_fd_sc_hd__buf_1 _11420_ (.A(_05376_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_2 _11421_ (.A0(_05499_),
    .A1(\core.cpuregs[30][16] ),
    .S(_05487_),
    .X(_05500_));
 sky130_fd_sc_hd__buf_1 _11422_ (.A(_05500_),
    .X(_00324_));
 sky130_fd_sc_hd__buf_1 _11423_ (.A(_05382_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_2 _11424_ (.A0(_05501_),
    .A1(\core.cpuregs[30][17] ),
    .S(_05487_),
    .X(_05502_));
 sky130_fd_sc_hd__buf_1 _11425_ (.A(_05502_),
    .X(_00325_));
 sky130_fd_sc_hd__buf_1 _11426_ (.A(_05387_),
    .X(_05503_));
 sky130_fd_sc_hd__mux2_2 _11427_ (.A0(_05503_),
    .A1(\core.cpuregs[30][18] ),
    .S(_05487_),
    .X(_05504_));
 sky130_fd_sc_hd__buf_1 _11428_ (.A(_05504_),
    .X(_00326_));
 sky130_fd_sc_hd__buf_1 _11429_ (.A(_05392_),
    .X(_05505_));
 sky130_fd_sc_hd__mux2_2 _11430_ (.A0(_05505_),
    .A1(\core.cpuregs[30][19] ),
    .S(_05487_),
    .X(_05506_));
 sky130_fd_sc_hd__buf_1 _11431_ (.A(_05506_),
    .X(_00327_));
 sky130_fd_sc_hd__buf_1 _11432_ (.A(_05398_),
    .X(_05507_));
 sky130_fd_sc_hd__buf_1 _11433_ (.A(_05465_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_2 _11434_ (.A0(_05507_),
    .A1(\core.cpuregs[30][20] ),
    .S(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__buf_1 _11435_ (.A(_05509_),
    .X(_00328_));
 sky130_fd_sc_hd__buf_1 _11436_ (.A(_05404_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_2 _11437_ (.A0(_05510_),
    .A1(\core.cpuregs[30][21] ),
    .S(_05508_),
    .X(_05511_));
 sky130_fd_sc_hd__buf_1 _11438_ (.A(_05511_),
    .X(_00329_));
 sky130_fd_sc_hd__buf_1 _11439_ (.A(_05409_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_2 _11440_ (.A0(_05512_),
    .A1(\core.cpuregs[30][22] ),
    .S(_05508_),
    .X(_05513_));
 sky130_fd_sc_hd__buf_1 _11441_ (.A(_05513_),
    .X(_00330_));
 sky130_fd_sc_hd__buf_1 _11442_ (.A(_05415_),
    .X(_05514_));
 sky130_fd_sc_hd__mux2_2 _11443_ (.A0(_05514_),
    .A1(\core.cpuregs[30][23] ),
    .S(_05508_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_1 _11444_ (.A(_05515_),
    .X(_00331_));
 sky130_fd_sc_hd__buf_1 _11445_ (.A(_05420_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_2 _11446_ (.A0(_05516_),
    .A1(\core.cpuregs[30][24] ),
    .S(_05508_),
    .X(_05517_));
 sky130_fd_sc_hd__buf_1 _11447_ (.A(_05517_),
    .X(_00332_));
 sky130_fd_sc_hd__buf_1 _11448_ (.A(_05425_),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_2 _11449_ (.A0(_05518_),
    .A1(\core.cpuregs[30][25] ),
    .S(_05508_),
    .X(_05519_));
 sky130_fd_sc_hd__buf_1 _11450_ (.A(_05519_),
    .X(_00333_));
 sky130_fd_sc_hd__buf_1 _11451_ (.A(_05431_),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_2 _11452_ (.A0(_05520_),
    .A1(\core.cpuregs[30][26] ),
    .S(_05508_),
    .X(_05521_));
 sky130_fd_sc_hd__buf_1 _11453_ (.A(_05521_),
    .X(_00334_));
 sky130_fd_sc_hd__buf_1 _11454_ (.A(_05436_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_2 _11455_ (.A0(_05522_),
    .A1(\core.cpuregs[30][27] ),
    .S(_05508_),
    .X(_05523_));
 sky130_fd_sc_hd__buf_1 _11456_ (.A(_05523_),
    .X(_00335_));
 sky130_fd_sc_hd__buf_1 _11457_ (.A(_05441_),
    .X(_05524_));
 sky130_fd_sc_hd__mux2_2 _11458_ (.A0(_05524_),
    .A1(\core.cpuregs[30][28] ),
    .S(_05508_),
    .X(_05525_));
 sky130_fd_sc_hd__buf_1 _11459_ (.A(_05525_),
    .X(_00336_));
 sky130_fd_sc_hd__buf_1 _11460_ (.A(_05447_),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_2 _11461_ (.A0(_05526_),
    .A1(\core.cpuregs[30][29] ),
    .S(_05508_),
    .X(_05527_));
 sky130_fd_sc_hd__buf_1 _11462_ (.A(_05527_),
    .X(_00337_));
 sky130_fd_sc_hd__buf_1 _11463_ (.A(_05452_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_2 _11464_ (.A0(_05528_),
    .A1(\core.cpuregs[30][30] ),
    .S(_05465_),
    .X(_05529_));
 sky130_fd_sc_hd__buf_1 _11465_ (.A(_05529_),
    .X(_00338_));
 sky130_fd_sc_hd__buf_1 _11466_ (.A(_05457_),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_2 _11467_ (.A0(_05530_),
    .A1(\core.cpuregs[30][31] ),
    .S(_05465_),
    .X(_05531_));
 sky130_fd_sc_hd__buf_1 _11468_ (.A(_05531_),
    .X(_00339_));
 sky130_fd_sc_hd__mux4_2 _11469_ (.A0(\core.cpuregs[4][0] ),
    .A1(\core.cpuregs[5][0] ),
    .A2(\core.cpuregs[6][0] ),
    .A3(\core.cpuregs[7][0] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_05532_));
 sky130_fd_sc_hd__or2_2 _11470_ (.A(_02132_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__mux4_2 _11471_ (.A0(\core.cpuregs[0][0] ),
    .A1(\core.cpuregs[1][0] ),
    .A2(\core.cpuregs[2][0] ),
    .A3(\core.cpuregs[3][0] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_05534_));
 sky130_fd_sc_hd__or2_2 _11472_ (.A(_02139_),
    .B(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__mux4_2 _11473_ (.A0(\core.cpuregs[8][0] ),
    .A1(\core.cpuregs[9][0] ),
    .A2(\core.cpuregs[10][0] ),
    .A3(\core.cpuregs[11][0] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_05536_));
 sky130_fd_sc_hd__or2_2 _11474_ (.A(_02139_),
    .B(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__mux4_2 _11475_ (.A0(\core.cpuregs[12][0] ),
    .A1(\core.cpuregs[13][0] ),
    .A2(\core.cpuregs[14][0] ),
    .A3(\core.cpuregs[15][0] ),
    .S0(_02149_),
    .S1(_02144_),
    .X(_05538_));
 sky130_fd_sc_hd__o21a_2 _11476_ (.A1(_02132_),
    .A2(_05538_),
    .B1(_02151_),
    .X(_05539_));
 sky130_fd_sc_hd__a32o_2 _11477_ (.A1(_02128_),
    .A2(_05533_),
    .A3(_05535_),
    .B1(_05537_),
    .B2(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__mux4_2 _11478_ (.A0(\core.cpuregs[24][0] ),
    .A1(\core.cpuregs[25][0] ),
    .A2(\core.cpuregs[26][0] ),
    .A3(\core.cpuregs[27][0] ),
    .S0(_02155_),
    .S1(_02156_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_2 _11479_ (.A0(\core.cpuregs[30][0] ),
    .A1(\core.cpuregs[31][0] ),
    .S(_02148_),
    .X(_05542_));
 sky130_fd_sc_hd__mux2_2 _11480_ (.A0(\core.cpuregs[28][0] ),
    .A1(\core.cpuregs[29][0] ),
    .S(_02133_),
    .X(_05543_));
 sky130_fd_sc_hd__a21o_2 _11481_ (.A1(_02161_),
    .A2(_05543_),
    .B1(_02131_),
    .X(_05544_));
 sky130_fd_sc_hd__a21o_2 _11482_ (.A1(_02144_),
    .A2(_05542_),
    .B1(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__o211a_2 _11483_ (.A1(_02138_),
    .A2(_05541_),
    .B1(_05545_),
    .C1(_02151_),
    .X(_05546_));
 sky130_fd_sc_hd__mux4_2 _11484_ (.A0(\core.cpuregs[20][0] ),
    .A1(\core.cpuregs[21][0] ),
    .A2(\core.cpuregs[22][0] ),
    .A3(\core.cpuregs[23][0] ),
    .S0(_02134_),
    .S1(_02156_),
    .X(_05547_));
 sky130_fd_sc_hd__mux2_2 _11485_ (.A0(\core.cpuregs[16][0] ),
    .A1(\core.cpuregs[17][0] ),
    .S(_02148_),
    .X(_05548_));
 sky130_fd_sc_hd__mux2_2 _11486_ (.A0(\core.cpuregs[18][0] ),
    .A1(\core.cpuregs[19][0] ),
    .S(_02133_),
    .X(_05549_));
 sky130_fd_sc_hd__a21o_2 _11487_ (.A1(_02158_),
    .A2(_05549_),
    .B1(_02138_),
    .X(_05550_));
 sky130_fd_sc_hd__a21o_2 _11488_ (.A1(_02161_),
    .A2(_05548_),
    .B1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o211a_2 _11489_ (.A1(_02131_),
    .A2(_05547_),
    .B1(_05551_),
    .C1(_02128_),
    .X(_05552_));
 sky130_fd_sc_hd__or3b_2 _11490_ (.A(_05546_),
    .B(_05552_),
    .C_N(_00004_),
    .X(_05553_));
 sky130_fd_sc_hd__o211a_2 _11491_ (.A1(_00004_),
    .A2(_05540_),
    .B1(_05553_),
    .C1(_02175_),
    .X(_05554_));
 sky130_fd_sc_hd__mux2_2 _11492_ (.A0(_05554_),
    .A1(\core.decoded_imm_j[11] ),
    .S(\core.is_slli_srli_srai ),
    .X(_05555_));
 sky130_fd_sc_hd__a21oi_2 _11493_ (.A1(\core.reg_sh[0] ),
    .A2(_02179_),
    .B1(_02126_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21o_2 _11494_ (.A1(_02126_),
    .A2(_05555_),
    .B1(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__o31a_2 _11495_ (.A1(_02126_),
    .A2(\core.reg_sh[0] ),
    .A3(_02179_),
    .B1(_05557_),
    .X(_00340_));
 sky130_fd_sc_hd__a21o_2 _11496_ (.A1(\core.reg_sh[0] ),
    .A2(\core.reg_sh[1] ),
    .B1(_02180_),
    .X(_05558_));
 sky130_fd_sc_hd__mux4_2 _11497_ (.A0(\core.cpuregs[4][1] ),
    .A1(\core.cpuregs[5][1] ),
    .A2(\core.cpuregs[6][1] ),
    .A3(\core.cpuregs[7][1] ),
    .S0(_02155_),
    .S1(_02158_),
    .X(_05559_));
 sky130_fd_sc_hd__or2_2 _11498_ (.A(_02131_),
    .B(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__mux4_2 _11499_ (.A0(\core.cpuregs[0][1] ),
    .A1(\core.cpuregs[1][1] ),
    .A2(\core.cpuregs[2][1] ),
    .A3(\core.cpuregs[3][1] ),
    .S0(_02155_),
    .S1(_02158_),
    .X(_05561_));
 sky130_fd_sc_hd__or2_2 _11500_ (.A(_02138_),
    .B(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__mux4_2 _11501_ (.A0(\core.cpuregs[8][1] ),
    .A1(\core.cpuregs[9][1] ),
    .A2(\core.cpuregs[10][1] ),
    .A3(\core.cpuregs[11][1] ),
    .S0(_02134_),
    .S1(_02135_),
    .X(_05563_));
 sky130_fd_sc_hd__or2_2 _11502_ (.A(_02139_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__mux4_2 _11503_ (.A0(\core.cpuregs[12][1] ),
    .A1(\core.cpuregs[13][1] ),
    .A2(\core.cpuregs[14][1] ),
    .A3(\core.cpuregs[15][1] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_05565_));
 sky130_fd_sc_hd__o21a_2 _11504_ (.A1(_02132_),
    .A2(_05565_),
    .B1(_02151_),
    .X(_05566_));
 sky130_fd_sc_hd__a32o_2 _11505_ (.A1(_02128_),
    .A2(_05560_),
    .A3(_05562_),
    .B1(_05564_),
    .B2(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__mux4_2 _11506_ (.A0(\core.cpuregs[24][1] ),
    .A1(\core.cpuregs[25][1] ),
    .A2(\core.cpuregs[26][1] ),
    .A3(\core.cpuregs[27][1] ),
    .S0(_02155_),
    .S1(_02158_),
    .X(_05568_));
 sky130_fd_sc_hd__mux2_2 _11507_ (.A0(\core.cpuregs[30][1] ),
    .A1(\core.cpuregs[31][1] ),
    .S(_02148_),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_2 _11508_ (.A0(\core.cpuregs[28][1] ),
    .A1(\core.cpuregs[29][1] ),
    .S(_00000_),
    .X(_05570_));
 sky130_fd_sc_hd__a21o_2 _11509_ (.A1(_02161_),
    .A2(_05570_),
    .B1(_02130_),
    .X(_05571_));
 sky130_fd_sc_hd__a21o_2 _11510_ (.A1(_02144_),
    .A2(_05569_),
    .B1(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__o211a_2 _11511_ (.A1(_02138_),
    .A2(_05568_),
    .B1(_05572_),
    .C1(_02151_),
    .X(_05573_));
 sky130_fd_sc_hd__mux4_2 _11512_ (.A0(\core.cpuregs[20][1] ),
    .A1(\core.cpuregs[21][1] ),
    .A2(\core.cpuregs[22][1] ),
    .A3(\core.cpuregs[23][1] ),
    .S0(_02155_),
    .S1(_02158_),
    .X(_05574_));
 sky130_fd_sc_hd__mux2_2 _11513_ (.A0(\core.cpuregs[16][1] ),
    .A1(\core.cpuregs[17][1] ),
    .S(_02148_),
    .X(_05575_));
 sky130_fd_sc_hd__mux2_2 _11514_ (.A0(\core.cpuregs[18][1] ),
    .A1(\core.cpuregs[19][1] ),
    .S(_00000_),
    .X(_05576_));
 sky130_fd_sc_hd__a21o_2 _11515_ (.A1(_02158_),
    .A2(_05576_),
    .B1(_00002_),
    .X(_05577_));
 sky130_fd_sc_hd__a21o_2 _11516_ (.A1(_02161_),
    .A2(_05575_),
    .B1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__o211a_2 _11517_ (.A1(_02131_),
    .A2(_05574_),
    .B1(_05578_),
    .C1(_02128_),
    .X(_05579_));
 sky130_fd_sc_hd__or3b_2 _11518_ (.A(_05573_),
    .B(_05579_),
    .C_N(_00004_),
    .X(_05580_));
 sky130_fd_sc_hd__o211a_2 _11519_ (.A1(_00004_),
    .A2(_05567_),
    .B1(_05580_),
    .C1(_02175_),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_2 _11520_ (.A0(_05581_),
    .A1(\core.decoded_imm_j[1] ),
    .S(\core.is_slli_srli_srai ),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_2 _11521_ (.A0(_05558_),
    .A1(_05582_),
    .S(_02126_),
    .X(_05583_));
 sky130_fd_sc_hd__o31a_2 _11522_ (.A1(_02126_),
    .A2(\core.reg_sh[1] ),
    .A3(_02179_),
    .B1(_05583_),
    .X(_00341_));
 sky130_fd_sc_hd__or2_2 _11523_ (.A(_05285_),
    .B(_05464_),
    .X(_05584_));
 sky130_fd_sc_hd__buf_1 _11524_ (.A(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_2 _11525_ (.A0(_05460_),
    .A1(\core.cpuregs[22][0] ),
    .S(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_1 _11526_ (.A(_05586_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_2 _11527_ (.A0(_05468_),
    .A1(\core.cpuregs[22][1] ),
    .S(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_1 _11528_ (.A(_05587_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_2 _11529_ (.A0(_05470_),
    .A1(\core.cpuregs[22][2] ),
    .S(_05585_),
    .X(_05588_));
 sky130_fd_sc_hd__buf_1 _11530_ (.A(_05588_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_2 _11531_ (.A0(_05472_),
    .A1(\core.cpuregs[22][3] ),
    .S(_05585_),
    .X(_05589_));
 sky130_fd_sc_hd__buf_1 _11532_ (.A(_05589_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_2 _11533_ (.A0(_05474_),
    .A1(\core.cpuregs[22][4] ),
    .S(_05585_),
    .X(_05590_));
 sky130_fd_sc_hd__buf_1 _11534_ (.A(_05590_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_2 _11535_ (.A0(_05476_),
    .A1(\core.cpuregs[22][5] ),
    .S(_05585_),
    .X(_05591_));
 sky130_fd_sc_hd__buf_1 _11536_ (.A(_05591_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_2 _11537_ (.A0(_05478_),
    .A1(\core.cpuregs[22][6] ),
    .S(_05585_),
    .X(_05592_));
 sky130_fd_sc_hd__buf_1 _11538_ (.A(_05592_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_2 _11539_ (.A0(_05480_),
    .A1(\core.cpuregs[22][7] ),
    .S(_05585_),
    .X(_05593_));
 sky130_fd_sc_hd__buf_1 _11540_ (.A(_05593_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_2 _11541_ (.A0(_05482_),
    .A1(\core.cpuregs[22][8] ),
    .S(_05585_),
    .X(_05594_));
 sky130_fd_sc_hd__buf_1 _11542_ (.A(_05594_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_2 _11543_ (.A0(_05484_),
    .A1(\core.cpuregs[22][9] ),
    .S(_05585_),
    .X(_05595_));
 sky130_fd_sc_hd__buf_1 _11544_ (.A(_05595_),
    .X(_00351_));
 sky130_fd_sc_hd__buf_1 _11545_ (.A(_05584_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_2 _11546_ (.A0(_05486_),
    .A1(\core.cpuregs[22][10] ),
    .S(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__buf_1 _11547_ (.A(_05597_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_2 _11548_ (.A0(_05489_),
    .A1(\core.cpuregs[22][11] ),
    .S(_05596_),
    .X(_05598_));
 sky130_fd_sc_hd__buf_1 _11549_ (.A(_05598_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_2 _11550_ (.A0(_05491_),
    .A1(\core.cpuregs[22][12] ),
    .S(_05596_),
    .X(_05599_));
 sky130_fd_sc_hd__buf_1 _11551_ (.A(_05599_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_2 _11552_ (.A0(_05493_),
    .A1(\core.cpuregs[22][13] ),
    .S(_05596_),
    .X(_05600_));
 sky130_fd_sc_hd__buf_1 _11553_ (.A(_05600_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_2 _11554_ (.A0(_05495_),
    .A1(\core.cpuregs[22][14] ),
    .S(_05596_),
    .X(_05601_));
 sky130_fd_sc_hd__buf_1 _11555_ (.A(_05601_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_2 _11556_ (.A0(_05497_),
    .A1(\core.cpuregs[22][15] ),
    .S(_05596_),
    .X(_05602_));
 sky130_fd_sc_hd__buf_1 _11557_ (.A(_05602_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_2 _11558_ (.A0(_05499_),
    .A1(\core.cpuregs[22][16] ),
    .S(_05596_),
    .X(_05603_));
 sky130_fd_sc_hd__buf_1 _11559_ (.A(_05603_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_2 _11560_ (.A0(_05501_),
    .A1(\core.cpuregs[22][17] ),
    .S(_05596_),
    .X(_05604_));
 sky130_fd_sc_hd__buf_1 _11561_ (.A(_05604_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_2 _11562_ (.A0(_05503_),
    .A1(\core.cpuregs[22][18] ),
    .S(_05596_),
    .X(_05605_));
 sky130_fd_sc_hd__buf_1 _11563_ (.A(_05605_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_2 _11564_ (.A0(_05505_),
    .A1(\core.cpuregs[22][19] ),
    .S(_05596_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_1 _11565_ (.A(_05606_),
    .X(_00361_));
 sky130_fd_sc_hd__buf_1 _11566_ (.A(_05584_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_2 _11567_ (.A0(_05507_),
    .A1(\core.cpuregs[22][20] ),
    .S(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__buf_1 _11568_ (.A(_05608_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_2 _11569_ (.A0(_05510_),
    .A1(\core.cpuregs[22][21] ),
    .S(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_1 _11570_ (.A(_05609_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_2 _11571_ (.A0(_05512_),
    .A1(\core.cpuregs[22][22] ),
    .S(_05607_),
    .X(_05610_));
 sky130_fd_sc_hd__buf_1 _11572_ (.A(_05610_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_2 _11573_ (.A0(_05514_),
    .A1(\core.cpuregs[22][23] ),
    .S(_05607_),
    .X(_05611_));
 sky130_fd_sc_hd__buf_1 _11574_ (.A(_05611_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_2 _11575_ (.A0(_05516_),
    .A1(\core.cpuregs[22][24] ),
    .S(_05607_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_1 _11576_ (.A(_05612_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_2 _11577_ (.A0(_05518_),
    .A1(\core.cpuregs[22][25] ),
    .S(_05607_),
    .X(_05613_));
 sky130_fd_sc_hd__buf_1 _11578_ (.A(_05613_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_2 _11579_ (.A0(_05520_),
    .A1(\core.cpuregs[22][26] ),
    .S(_05607_),
    .X(_05614_));
 sky130_fd_sc_hd__buf_1 _11580_ (.A(_05614_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_2 _11581_ (.A0(_05522_),
    .A1(\core.cpuregs[22][27] ),
    .S(_05607_),
    .X(_05615_));
 sky130_fd_sc_hd__buf_1 _11582_ (.A(_05615_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_2 _11583_ (.A0(_05524_),
    .A1(\core.cpuregs[22][28] ),
    .S(_05607_),
    .X(_05616_));
 sky130_fd_sc_hd__buf_1 _11584_ (.A(_05616_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_2 _11585_ (.A0(_05526_),
    .A1(\core.cpuregs[22][29] ),
    .S(_05607_),
    .X(_05617_));
 sky130_fd_sc_hd__buf_1 _11586_ (.A(_05617_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_2 _11587_ (.A0(_05528_),
    .A1(\core.cpuregs[22][30] ),
    .S(_05584_),
    .X(_05618_));
 sky130_fd_sc_hd__buf_1 _11588_ (.A(_05618_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_2 _11589_ (.A0(_05530_),
    .A1(\core.cpuregs[22][31] ),
    .S(_05584_),
    .X(_05619_));
 sky130_fd_sc_hd__buf_1 _11590_ (.A(_05619_),
    .X(_00373_));
 sky130_fd_sc_hd__or3_2 _11591_ (.A(\core.latched_rd[4] ),
    .B(\core.latched_rd[3] ),
    .C(\core.latched_rd[2] ),
    .X(_05620_));
 sky130_fd_sc_hd__or2_2 _11592_ (.A(_05464_),
    .B(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__buf_1 _11593_ (.A(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__mux2_2 _11594_ (.A0(_05460_),
    .A1(\core.cpuregs[2][0] ),
    .S(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__buf_1 _11595_ (.A(_05623_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_2 _11596_ (.A0(_05468_),
    .A1(\core.cpuregs[2][1] ),
    .S(_05622_),
    .X(_05624_));
 sky130_fd_sc_hd__buf_1 _11597_ (.A(_05624_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_2 _11598_ (.A0(_05470_),
    .A1(\core.cpuregs[2][2] ),
    .S(_05622_),
    .X(_05625_));
 sky130_fd_sc_hd__buf_1 _11599_ (.A(_05625_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_2 _11600_ (.A0(_05472_),
    .A1(\core.cpuregs[2][3] ),
    .S(_05622_),
    .X(_05626_));
 sky130_fd_sc_hd__buf_1 _11601_ (.A(_05626_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_2 _11602_ (.A0(_05474_),
    .A1(\core.cpuregs[2][4] ),
    .S(_05622_),
    .X(_05627_));
 sky130_fd_sc_hd__buf_1 _11603_ (.A(_05627_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_2 _11604_ (.A0(_05476_),
    .A1(\core.cpuregs[2][5] ),
    .S(_05622_),
    .X(_05628_));
 sky130_fd_sc_hd__buf_1 _11605_ (.A(_05628_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_2 _11606_ (.A0(_05478_),
    .A1(\core.cpuregs[2][6] ),
    .S(_05622_),
    .X(_05629_));
 sky130_fd_sc_hd__buf_1 _11607_ (.A(_05629_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_2 _11608_ (.A0(_05480_),
    .A1(\core.cpuregs[2][7] ),
    .S(_05622_),
    .X(_05630_));
 sky130_fd_sc_hd__buf_1 _11609_ (.A(_05630_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_2 _11610_ (.A0(_05482_),
    .A1(\core.cpuregs[2][8] ),
    .S(_05622_),
    .X(_05631_));
 sky130_fd_sc_hd__buf_1 _11611_ (.A(_05631_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_2 _11612_ (.A0(_05484_),
    .A1(\core.cpuregs[2][9] ),
    .S(_05622_),
    .X(_05632_));
 sky130_fd_sc_hd__buf_1 _11613_ (.A(_05632_),
    .X(_00383_));
 sky130_fd_sc_hd__buf_1 _11614_ (.A(_05621_),
    .X(_05633_));
 sky130_fd_sc_hd__mux2_2 _11615_ (.A0(_05486_),
    .A1(\core.cpuregs[2][10] ),
    .S(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__buf_1 _11616_ (.A(_05634_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_2 _11617_ (.A0(_05489_),
    .A1(\core.cpuregs[2][11] ),
    .S(_05633_),
    .X(_05635_));
 sky130_fd_sc_hd__buf_1 _11618_ (.A(_05635_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_2 _11619_ (.A0(_05491_),
    .A1(\core.cpuregs[2][12] ),
    .S(_05633_),
    .X(_05636_));
 sky130_fd_sc_hd__buf_1 _11620_ (.A(_05636_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_2 _11621_ (.A0(_05493_),
    .A1(\core.cpuregs[2][13] ),
    .S(_05633_),
    .X(_05637_));
 sky130_fd_sc_hd__buf_1 _11622_ (.A(_05637_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_2 _11623_ (.A0(_05495_),
    .A1(\core.cpuregs[2][14] ),
    .S(_05633_),
    .X(_05638_));
 sky130_fd_sc_hd__buf_1 _11624_ (.A(_05638_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_2 _11625_ (.A0(_05497_),
    .A1(\core.cpuregs[2][15] ),
    .S(_05633_),
    .X(_05639_));
 sky130_fd_sc_hd__buf_1 _11626_ (.A(_05639_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_2 _11627_ (.A0(_05499_),
    .A1(\core.cpuregs[2][16] ),
    .S(_05633_),
    .X(_05640_));
 sky130_fd_sc_hd__buf_1 _11628_ (.A(_05640_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_2 _11629_ (.A0(_05501_),
    .A1(\core.cpuregs[2][17] ),
    .S(_05633_),
    .X(_05641_));
 sky130_fd_sc_hd__buf_1 _11630_ (.A(_05641_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_2 _11631_ (.A0(_05503_),
    .A1(\core.cpuregs[2][18] ),
    .S(_05633_),
    .X(_05642_));
 sky130_fd_sc_hd__buf_1 _11632_ (.A(_05642_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_2 _11633_ (.A0(_05505_),
    .A1(\core.cpuregs[2][19] ),
    .S(_05633_),
    .X(_05643_));
 sky130_fd_sc_hd__buf_1 _11634_ (.A(_05643_),
    .X(_00393_));
 sky130_fd_sc_hd__buf_1 _11635_ (.A(_05621_),
    .X(_05644_));
 sky130_fd_sc_hd__mux2_2 _11636_ (.A0(_05507_),
    .A1(\core.cpuregs[2][20] ),
    .S(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__buf_1 _11637_ (.A(_05645_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_2 _11638_ (.A0(_05510_),
    .A1(\core.cpuregs[2][21] ),
    .S(_05644_),
    .X(_05646_));
 sky130_fd_sc_hd__buf_1 _11639_ (.A(_05646_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_2 _11640_ (.A0(_05512_),
    .A1(\core.cpuregs[2][22] ),
    .S(_05644_),
    .X(_05647_));
 sky130_fd_sc_hd__buf_1 _11641_ (.A(_05647_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_2 _11642_ (.A0(_05514_),
    .A1(\core.cpuregs[2][23] ),
    .S(_05644_),
    .X(_05648_));
 sky130_fd_sc_hd__buf_1 _11643_ (.A(_05648_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_2 _11644_ (.A0(_05516_),
    .A1(\core.cpuregs[2][24] ),
    .S(_05644_),
    .X(_05649_));
 sky130_fd_sc_hd__buf_1 _11645_ (.A(_05649_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_2 _11646_ (.A0(_05518_),
    .A1(\core.cpuregs[2][25] ),
    .S(_05644_),
    .X(_05650_));
 sky130_fd_sc_hd__buf_1 _11647_ (.A(_05650_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_2 _11648_ (.A0(_05520_),
    .A1(\core.cpuregs[2][26] ),
    .S(_05644_),
    .X(_05651_));
 sky130_fd_sc_hd__buf_1 _11649_ (.A(_05651_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_2 _11650_ (.A0(_05522_),
    .A1(\core.cpuregs[2][27] ),
    .S(_05644_),
    .X(_05652_));
 sky130_fd_sc_hd__buf_1 _11651_ (.A(_05652_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_2 _11652_ (.A0(_05524_),
    .A1(\core.cpuregs[2][28] ),
    .S(_05644_),
    .X(_05653_));
 sky130_fd_sc_hd__buf_1 _11653_ (.A(_05653_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_2 _11654_ (.A0(_05526_),
    .A1(\core.cpuregs[2][29] ),
    .S(_05644_),
    .X(_05654_));
 sky130_fd_sc_hd__buf_1 _11655_ (.A(_05654_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_2 _11656_ (.A0(_05528_),
    .A1(\core.cpuregs[2][30] ),
    .S(_05621_),
    .X(_05655_));
 sky130_fd_sc_hd__buf_1 _11657_ (.A(_05655_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_2 _11658_ (.A0(_05530_),
    .A1(\core.cpuregs[2][31] ),
    .S(_05621_),
    .X(_05656_));
 sky130_fd_sc_hd__buf_1 _11659_ (.A(_05656_),
    .X(_00405_));
 sky130_fd_sc_hd__nand3b_2 _11660_ (.A_N(\core.latched_rd[2] ),
    .B(\core.latched_rd[3] ),
    .C(\core.latched_rd[4] ),
    .Y(_05657_));
 sky130_fd_sc_hd__nor2_2 _11661_ (.A(_05286_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__buf_1 _11662_ (.A(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_2 _11663_ (.A0(\core.cpuregs[27][0] ),
    .A1(_05284_),
    .S(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__buf_1 _11664_ (.A(_05660_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_2 _11665_ (.A0(\core.cpuregs[27][1] ),
    .A1(_05292_),
    .S(_05659_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _11666_ (.A(_05661_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_2 _11667_ (.A0(\core.cpuregs[27][2] ),
    .A1(_05297_),
    .S(_05659_),
    .X(_05662_));
 sky130_fd_sc_hd__buf_1 _11668_ (.A(_05662_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_2 _11669_ (.A0(\core.cpuregs[27][3] ),
    .A1(_05304_),
    .S(_05659_),
    .X(_05663_));
 sky130_fd_sc_hd__buf_1 _11670_ (.A(_05663_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_2 _11671_ (.A0(\core.cpuregs[27][4] ),
    .A1(_05310_),
    .S(_05659_),
    .X(_05664_));
 sky130_fd_sc_hd__buf_1 _11672_ (.A(_05664_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_2 _11673_ (.A0(\core.cpuregs[27][5] ),
    .A1(_05315_),
    .S(_05659_),
    .X(_05665_));
 sky130_fd_sc_hd__buf_1 _11674_ (.A(_05665_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_2 _11675_ (.A0(\core.cpuregs[27][6] ),
    .A1(_05320_),
    .S(_05659_),
    .X(_05666_));
 sky130_fd_sc_hd__buf_1 _11676_ (.A(_05666_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_2 _11677_ (.A0(\core.cpuregs[27][7] ),
    .A1(_05326_),
    .S(_05659_),
    .X(_05667_));
 sky130_fd_sc_hd__buf_1 _11678_ (.A(_05667_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_2 _11679_ (.A0(\core.cpuregs[27][8] ),
    .A1(_05332_),
    .S(_05659_),
    .X(_05668_));
 sky130_fd_sc_hd__buf_1 _11680_ (.A(_05668_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_2 _11681_ (.A0(\core.cpuregs[27][9] ),
    .A1(_05337_),
    .S(_05659_),
    .X(_05669_));
 sky130_fd_sc_hd__buf_1 _11682_ (.A(_05669_),
    .X(_00415_));
 sky130_fd_sc_hd__buf_1 _11683_ (.A(_05658_),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_2 _11684_ (.A0(\core.cpuregs[27][10] ),
    .A1(_05343_),
    .S(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__buf_1 _11685_ (.A(_05671_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_2 _11686_ (.A0(\core.cpuregs[27][11] ),
    .A1(_05349_),
    .S(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__buf_1 _11687_ (.A(_05672_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_2 _11688_ (.A0(\core.cpuregs[27][12] ),
    .A1(_05355_),
    .S(_05670_),
    .X(_05673_));
 sky130_fd_sc_hd__buf_1 _11689_ (.A(_05673_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_2 _11690_ (.A0(\core.cpuregs[27][13] ),
    .A1(_05360_),
    .S(_05670_),
    .X(_05674_));
 sky130_fd_sc_hd__buf_1 _11691_ (.A(_05674_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_2 _11692_ (.A0(\core.cpuregs[27][14] ),
    .A1(_05367_),
    .S(_05670_),
    .X(_05675_));
 sky130_fd_sc_hd__buf_1 _11693_ (.A(_05675_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_2 _11694_ (.A0(\core.cpuregs[27][15] ),
    .A1(_05372_),
    .S(_05670_),
    .X(_05676_));
 sky130_fd_sc_hd__buf_1 _11695_ (.A(_05676_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_2 _11696_ (.A0(\core.cpuregs[27][16] ),
    .A1(_05377_),
    .S(_05670_),
    .X(_05677_));
 sky130_fd_sc_hd__buf_1 _11697_ (.A(_05677_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_2 _11698_ (.A0(\core.cpuregs[27][17] ),
    .A1(_05383_),
    .S(_05670_),
    .X(_05678_));
 sky130_fd_sc_hd__buf_1 _11699_ (.A(_05678_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_2 _11700_ (.A0(\core.cpuregs[27][18] ),
    .A1(_05388_),
    .S(_05670_),
    .X(_05679_));
 sky130_fd_sc_hd__buf_1 _11701_ (.A(_05679_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_2 _11702_ (.A0(\core.cpuregs[27][19] ),
    .A1(_05393_),
    .S(_05670_),
    .X(_05680_));
 sky130_fd_sc_hd__buf_1 _11703_ (.A(_05680_),
    .X(_00425_));
 sky130_fd_sc_hd__buf_1 _11704_ (.A(_05658_),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_2 _11705_ (.A0(\core.cpuregs[27][20] ),
    .A1(_05399_),
    .S(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__buf_1 _11706_ (.A(_05682_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_2 _11707_ (.A0(\core.cpuregs[27][21] ),
    .A1(_05405_),
    .S(_05681_),
    .X(_05683_));
 sky130_fd_sc_hd__buf_1 _11708_ (.A(_05683_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_2 _11709_ (.A0(\core.cpuregs[27][22] ),
    .A1(_05410_),
    .S(_05681_),
    .X(_05684_));
 sky130_fd_sc_hd__buf_1 _11710_ (.A(_05684_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_2 _11711_ (.A0(\core.cpuregs[27][23] ),
    .A1(_05416_),
    .S(_05681_),
    .X(_05685_));
 sky130_fd_sc_hd__buf_1 _11712_ (.A(_05685_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_2 _11713_ (.A0(\core.cpuregs[27][24] ),
    .A1(_05421_),
    .S(_05681_),
    .X(_05686_));
 sky130_fd_sc_hd__buf_1 _11714_ (.A(_05686_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_2 _11715_ (.A0(\core.cpuregs[27][25] ),
    .A1(_05426_),
    .S(_05681_),
    .X(_05687_));
 sky130_fd_sc_hd__buf_1 _11716_ (.A(_05687_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_2 _11717_ (.A0(\core.cpuregs[27][26] ),
    .A1(_05432_),
    .S(_05681_),
    .X(_05688_));
 sky130_fd_sc_hd__buf_1 _11718_ (.A(_05688_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_2 _11719_ (.A0(\core.cpuregs[27][27] ),
    .A1(_05437_),
    .S(_05681_),
    .X(_05689_));
 sky130_fd_sc_hd__buf_1 _11720_ (.A(_05689_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_2 _11721_ (.A0(\core.cpuregs[27][28] ),
    .A1(_05442_),
    .S(_05681_),
    .X(_05690_));
 sky130_fd_sc_hd__buf_1 _11722_ (.A(_05690_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_2 _11723_ (.A0(\core.cpuregs[27][29] ),
    .A1(_05448_),
    .S(_05681_),
    .X(_05691_));
 sky130_fd_sc_hd__buf_1 _11724_ (.A(_05691_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_2 _11725_ (.A0(\core.cpuregs[27][30] ),
    .A1(_05453_),
    .S(_05658_),
    .X(_05692_));
 sky130_fd_sc_hd__buf_1 _11726_ (.A(_05692_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_2 _11727_ (.A0(\core.cpuregs[27][31] ),
    .A1(_05458_),
    .S(_05658_),
    .X(_05693_));
 sky130_fd_sc_hd__buf_1 _11728_ (.A(_05693_),
    .X(_00437_));
 sky130_fd_sc_hd__nor2_2 _11729_ (.A(_03211_),
    .B(_05269_),
    .Y(_05694_));
 sky130_fd_sc_hd__buf_1 _11730_ (.A(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__mux2_2 _11731_ (.A0(mem_wdata[0]),
    .A1(_02368_),
    .S(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__buf_1 _11732_ (.A(_05696_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_2 _11733_ (.A0(mem_wdata[1]),
    .A1(_02366_),
    .S(_05695_),
    .X(_05697_));
 sky130_fd_sc_hd__buf_1 _11734_ (.A(_05697_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_2 _11735_ (.A0(mem_wdata[2]),
    .A1(\core.mem_la_wdata[2] ),
    .S(_05695_),
    .X(_05698_));
 sky130_fd_sc_hd__buf_1 _11736_ (.A(_05698_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_2 _11737_ (.A0(mem_wdata[3]),
    .A1(\core.mem_la_wdata[3] ),
    .S(_05695_),
    .X(_05699_));
 sky130_fd_sc_hd__buf_1 _11738_ (.A(_05699_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_2 _11739_ (.A0(mem_wdata[4]),
    .A1(\core.mem_la_wdata[4] ),
    .S(_05695_),
    .X(_05700_));
 sky130_fd_sc_hd__buf_1 _11740_ (.A(_05700_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_2 _11741_ (.A0(mem_wdata[5]),
    .A1(\core.mem_la_wdata[5] ),
    .S(_05695_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_1 _11742_ (.A(_05701_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_2 _11743_ (.A0(mem_wdata[6]),
    .A1(\core.mem_la_wdata[6] ),
    .S(_05695_),
    .X(_05702_));
 sky130_fd_sc_hd__buf_1 _11744_ (.A(_05702_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_2 _11745_ (.A0(mem_wdata[7]),
    .A1(\core.mem_la_wdata[7] ),
    .S(_05695_),
    .X(_05703_));
 sky130_fd_sc_hd__buf_1 _11746_ (.A(_05703_),
    .X(_00445_));
 sky130_fd_sc_hd__buf_1 _11747_ (.A(_02695_),
    .X(_05704_));
 sky130_fd_sc_hd__a22o_2 _11748_ (.A1(_02023_),
    .A2(_02368_),
    .B1(\core.pcpi_rs2[8] ),
    .B2(_02123_),
    .X(_05705_));
 sky130_fd_sc_hd__a21o_2 _11749_ (.A1(\core.pcpi_rs2[8] ),
    .A2(_05704_),
    .B1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__mux2_2 _11750_ (.A0(mem_wdata[8]),
    .A1(_05706_),
    .S(_05695_),
    .X(_05707_));
 sky130_fd_sc_hd__buf_1 _11751_ (.A(_05707_),
    .X(_00446_));
 sky130_fd_sc_hd__a22o_2 _11752_ (.A1(_02023_),
    .A2(_02366_),
    .B1(\core.pcpi_rs2[9] ),
    .B2(_02123_),
    .X(_05708_));
 sky130_fd_sc_hd__a21o_2 _11753_ (.A1(\core.pcpi_rs2[9] ),
    .A2(_05704_),
    .B1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__mux2_2 _11754_ (.A0(mem_wdata[9]),
    .A1(_05709_),
    .S(_05695_),
    .X(_05710_));
 sky130_fd_sc_hd__buf_1 _11755_ (.A(_05710_),
    .X(_00447_));
 sky130_fd_sc_hd__a22o_2 _11756_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[2] ),
    .B1(\core.pcpi_rs2[10] ),
    .B2(_02123_),
    .X(_05711_));
 sky130_fd_sc_hd__a21o_2 _11757_ (.A1(\core.pcpi_rs2[10] ),
    .A2(_05704_),
    .B1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _11758_ (.A(_05694_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_2 _11759_ (.A0(mem_wdata[10]),
    .A1(_05712_),
    .S(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__buf_1 _11760_ (.A(_05714_),
    .X(_00448_));
 sky130_fd_sc_hd__a22o_2 _11761_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[3] ),
    .B1(\core.pcpi_rs2[11] ),
    .B2(_02123_),
    .X(_05715_));
 sky130_fd_sc_hd__a21o_2 _11762_ (.A1(\core.pcpi_rs2[11] ),
    .A2(_05704_),
    .B1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_2 _11763_ (.A0(mem_wdata[11]),
    .A1(_05716_),
    .S(_05713_),
    .X(_05717_));
 sky130_fd_sc_hd__buf_1 _11764_ (.A(_05717_),
    .X(_00449_));
 sky130_fd_sc_hd__a22o_2 _11765_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[4] ),
    .B1(\core.pcpi_rs2[12] ),
    .B2(_02069_),
    .X(_05718_));
 sky130_fd_sc_hd__a21o_2 _11766_ (.A1(\core.pcpi_rs2[12] ),
    .A2(_05704_),
    .B1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__mux2_2 _11767_ (.A0(mem_wdata[12]),
    .A1(_05719_),
    .S(_05713_),
    .X(_05720_));
 sky130_fd_sc_hd__buf_1 _11768_ (.A(_05720_),
    .X(_00450_));
 sky130_fd_sc_hd__a22o_2 _11769_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[5] ),
    .B1(\core.pcpi_rs2[13] ),
    .B2(_02069_),
    .X(_05721_));
 sky130_fd_sc_hd__a21o_2 _11770_ (.A1(\core.pcpi_rs2[13] ),
    .A2(_05704_),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__mux2_2 _11771_ (.A0(mem_wdata[13]),
    .A1(_05722_),
    .S(_05713_),
    .X(_05723_));
 sky130_fd_sc_hd__buf_1 _11772_ (.A(_05723_),
    .X(_00451_));
 sky130_fd_sc_hd__a22o_2 _11773_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[6] ),
    .B1(\core.pcpi_rs2[14] ),
    .B2(_02069_),
    .X(_05724_));
 sky130_fd_sc_hd__a21o_2 _11774_ (.A1(\core.pcpi_rs2[14] ),
    .A2(_05704_),
    .B1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__mux2_2 _11775_ (.A0(mem_wdata[14]),
    .A1(_05725_),
    .S(_05713_),
    .X(_05726_));
 sky130_fd_sc_hd__buf_1 _11776_ (.A(_05726_),
    .X(_00452_));
 sky130_fd_sc_hd__a22o_2 _11777_ (.A1(_02023_),
    .A2(\core.mem_la_wdata[7] ),
    .B1(\core.pcpi_rs2[15] ),
    .B2(_02069_),
    .X(_05727_));
 sky130_fd_sc_hd__a21o_2 _11778_ (.A1(\core.pcpi_rs2[15] ),
    .A2(_05704_),
    .B1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_2 _11779_ (.A0(mem_wdata[15]),
    .A1(_05728_),
    .S(_05713_),
    .X(_05729_));
 sky130_fd_sc_hd__buf_1 _11780_ (.A(_05729_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_2 _11781_ (.A0(_02368_),
    .A1(\core.pcpi_rs2[16] ),
    .S(_02722_),
    .X(_05730_));
 sky130_fd_sc_hd__mux2_2 _11782_ (.A0(mem_wdata[16]),
    .A1(_05730_),
    .S(_05713_),
    .X(_05731_));
 sky130_fd_sc_hd__buf_1 _11783_ (.A(_05731_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_2 _11784_ (.A0(_02366_),
    .A1(\core.pcpi_rs2[17] ),
    .S(_02722_),
    .X(_05732_));
 sky130_fd_sc_hd__mux2_2 _11785_ (.A0(mem_wdata[17]),
    .A1(_05732_),
    .S(_05713_),
    .X(_05733_));
 sky130_fd_sc_hd__buf_1 _11786_ (.A(_05733_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_2 _11787_ (.A0(\core.mem_la_wdata[2] ),
    .A1(\core.pcpi_rs2[18] ),
    .S(_02722_),
    .X(_05734_));
 sky130_fd_sc_hd__mux2_2 _11788_ (.A0(mem_wdata[18]),
    .A1(_05734_),
    .S(_05713_),
    .X(_05735_));
 sky130_fd_sc_hd__buf_1 _11789_ (.A(_05735_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_2 _11790_ (.A0(\core.mem_la_wdata[3] ),
    .A1(\core.pcpi_rs2[19] ),
    .S(_02722_),
    .X(_05736_));
 sky130_fd_sc_hd__mux2_2 _11791_ (.A0(mem_wdata[19]),
    .A1(_05736_),
    .S(_05713_),
    .X(_05737_));
 sky130_fd_sc_hd__buf_1 _11792_ (.A(_05737_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_2 _11793_ (.A0(\core.mem_la_wdata[4] ),
    .A1(\core.pcpi_rs2[20] ),
    .S(_02695_),
    .X(_05738_));
 sky130_fd_sc_hd__buf_1 _11794_ (.A(_05694_),
    .X(_05739_));
 sky130_fd_sc_hd__mux2_2 _11795_ (.A0(mem_wdata[20]),
    .A1(_05738_),
    .S(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__buf_1 _11796_ (.A(_05740_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_2 _11797_ (.A0(\core.mem_la_wdata[5] ),
    .A1(\core.pcpi_rs2[21] ),
    .S(_02695_),
    .X(_05741_));
 sky130_fd_sc_hd__mux2_2 _11798_ (.A0(mem_wdata[21]),
    .A1(_05741_),
    .S(_05739_),
    .X(_05742_));
 sky130_fd_sc_hd__buf_1 _11799_ (.A(_05742_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_2 _11800_ (.A0(\core.mem_la_wdata[6] ),
    .A1(\core.pcpi_rs2[22] ),
    .S(_02695_),
    .X(_05743_));
 sky130_fd_sc_hd__mux2_2 _11801_ (.A0(mem_wdata[22]),
    .A1(_05743_),
    .S(_05739_),
    .X(_05744_));
 sky130_fd_sc_hd__buf_1 _11802_ (.A(_05744_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_2 _11803_ (.A0(\core.mem_la_wdata[7] ),
    .A1(\core.pcpi_rs2[23] ),
    .S(_02695_),
    .X(_05745_));
 sky130_fd_sc_hd__mux2_2 _11804_ (.A0(mem_wdata[23]),
    .A1(_05745_),
    .S(_05739_),
    .X(_05746_));
 sky130_fd_sc_hd__buf_1 _11805_ (.A(_05746_),
    .X(_00461_));
 sky130_fd_sc_hd__a21o_2 _11806_ (.A1(\core.pcpi_rs2[24] ),
    .A2(_05704_),
    .B1(_05705_),
    .X(_05747_));
 sky130_fd_sc_hd__mux2_2 _11807_ (.A0(mem_wdata[24]),
    .A1(_05747_),
    .S(_05739_),
    .X(_05748_));
 sky130_fd_sc_hd__buf_1 _11808_ (.A(_05748_),
    .X(_00462_));
 sky130_fd_sc_hd__a21o_2 _11809_ (.A1(\core.pcpi_rs2[25] ),
    .A2(_02708_),
    .B1(_05708_),
    .X(_05749_));
 sky130_fd_sc_hd__mux2_2 _11810_ (.A0(mem_wdata[25]),
    .A1(_05749_),
    .S(_05739_),
    .X(_05750_));
 sky130_fd_sc_hd__buf_1 _11811_ (.A(_05750_),
    .X(_00463_));
 sky130_fd_sc_hd__a21o_2 _11812_ (.A1(\core.pcpi_rs2[26] ),
    .A2(_02708_),
    .B1(_05711_),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_2 _11813_ (.A0(mem_wdata[26]),
    .A1(_05751_),
    .S(_05739_),
    .X(_05752_));
 sky130_fd_sc_hd__buf_1 _11814_ (.A(_05752_),
    .X(_00464_));
 sky130_fd_sc_hd__a21o_2 _11815_ (.A1(\core.pcpi_rs2[27] ),
    .A2(_02708_),
    .B1(_05715_),
    .X(_05753_));
 sky130_fd_sc_hd__mux2_2 _11816_ (.A0(mem_wdata[27]),
    .A1(_05753_),
    .S(_05739_),
    .X(_05754_));
 sky130_fd_sc_hd__buf_1 _11817_ (.A(_05754_),
    .X(_00465_));
 sky130_fd_sc_hd__a21o_2 _11818_ (.A1(\core.pcpi_rs2[28] ),
    .A2(_02708_),
    .B1(_05718_),
    .X(_05755_));
 sky130_fd_sc_hd__mux2_2 _11819_ (.A0(mem_wdata[28]),
    .A1(_05755_),
    .S(_05739_),
    .X(_05756_));
 sky130_fd_sc_hd__buf_1 _11820_ (.A(_05756_),
    .X(_00466_));
 sky130_fd_sc_hd__a21o_2 _11821_ (.A1(\core.pcpi_rs2[29] ),
    .A2(_02708_),
    .B1(_05721_),
    .X(_05757_));
 sky130_fd_sc_hd__mux2_2 _11822_ (.A0(mem_wdata[29]),
    .A1(_05757_),
    .S(_05739_),
    .X(_05758_));
 sky130_fd_sc_hd__buf_1 _11823_ (.A(_05758_),
    .X(_00467_));
 sky130_fd_sc_hd__a21o_2 _11824_ (.A1(\core.pcpi_rs2[30] ),
    .A2(_02708_),
    .B1(_05724_),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_2 _11825_ (.A0(mem_wdata[30]),
    .A1(_05759_),
    .S(_05694_),
    .X(_05760_));
 sky130_fd_sc_hd__buf_1 _11826_ (.A(_05760_),
    .X(_00468_));
 sky130_fd_sc_hd__a21o_2 _11827_ (.A1(\core.pcpi_rs2[31] ),
    .A2(_02708_),
    .B1(_05727_),
    .X(_05761_));
 sky130_fd_sc_hd__mux2_2 _11828_ (.A0(mem_wdata[31]),
    .A1(_05761_),
    .S(_05694_),
    .X(_05762_));
 sky130_fd_sc_hd__buf_1 _11829_ (.A(_05762_),
    .X(_00469_));
 sky130_fd_sc_hd__and2b_2 _11830_ (.A_N(\core.mem_do_wdata ),
    .B(_03207_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_2 _11831_ (.A0(mem_instr),
    .A1(_05763_),
    .S(_03236_),
    .X(_05764_));
 sky130_fd_sc_hd__buf_1 _11832_ (.A(_05764_),
    .X(_00470_));
 sky130_fd_sc_hd__or4b_2 _11833_ (.A(\core.latched_rd[1] ),
    .B(\core.latched_rd[0] ),
    .C(_05462_),
    .D_N(_05620_),
    .X(_05765_));
 sky130_fd_sc_hd__buf_1 _11834_ (.A(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__nor2_2 _11835_ (.A(_05461_),
    .B(_05766_),
    .Y(_05767_));
 sky130_fd_sc_hd__buf_1 _11836_ (.A(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__mux2_2 _11837_ (.A0(\core.cpuregs[28][0] ),
    .A1(_05284_),
    .S(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__buf_1 _11838_ (.A(_05769_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_2 _11839_ (.A0(\core.cpuregs[28][1] ),
    .A1(_05292_),
    .S(_05768_),
    .X(_05770_));
 sky130_fd_sc_hd__buf_1 _11840_ (.A(_05770_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_2 _11841_ (.A0(\core.cpuregs[28][2] ),
    .A1(_05297_),
    .S(_05768_),
    .X(_05771_));
 sky130_fd_sc_hd__buf_1 _11842_ (.A(_05771_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_2 _11843_ (.A0(\core.cpuregs[28][3] ),
    .A1(_05304_),
    .S(_05768_),
    .X(_05772_));
 sky130_fd_sc_hd__buf_1 _11844_ (.A(_05772_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_2 _11845_ (.A0(\core.cpuregs[28][4] ),
    .A1(_05310_),
    .S(_05768_),
    .X(_05773_));
 sky130_fd_sc_hd__buf_1 _11846_ (.A(_05773_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_2 _11847_ (.A0(\core.cpuregs[28][5] ),
    .A1(_05315_),
    .S(_05768_),
    .X(_05774_));
 sky130_fd_sc_hd__buf_1 _11848_ (.A(_05774_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_2 _11849_ (.A0(\core.cpuregs[28][6] ),
    .A1(_05320_),
    .S(_05768_),
    .X(_05775_));
 sky130_fd_sc_hd__buf_1 _11850_ (.A(_05775_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_2 _11851_ (.A0(\core.cpuregs[28][7] ),
    .A1(_05326_),
    .S(_05768_),
    .X(_05776_));
 sky130_fd_sc_hd__buf_1 _11852_ (.A(_05776_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_2 _11853_ (.A0(\core.cpuregs[28][8] ),
    .A1(_05332_),
    .S(_05768_),
    .X(_05777_));
 sky130_fd_sc_hd__buf_1 _11854_ (.A(_05777_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_2 _11855_ (.A0(\core.cpuregs[28][9] ),
    .A1(_05337_),
    .S(_05768_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_1 _11856_ (.A(_05778_),
    .X(_00480_));
 sky130_fd_sc_hd__buf_1 _11857_ (.A(_05767_),
    .X(_05779_));
 sky130_fd_sc_hd__mux2_2 _11858_ (.A0(\core.cpuregs[28][10] ),
    .A1(_05343_),
    .S(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__buf_1 _11859_ (.A(_05780_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_2 _11860_ (.A0(\core.cpuregs[28][11] ),
    .A1(_05349_),
    .S(_05779_),
    .X(_05781_));
 sky130_fd_sc_hd__buf_1 _11861_ (.A(_05781_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_2 _11862_ (.A0(\core.cpuregs[28][12] ),
    .A1(_05355_),
    .S(_05779_),
    .X(_05782_));
 sky130_fd_sc_hd__buf_1 _11863_ (.A(_05782_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_2 _11864_ (.A0(\core.cpuregs[28][13] ),
    .A1(_05360_),
    .S(_05779_),
    .X(_05783_));
 sky130_fd_sc_hd__buf_1 _11865_ (.A(_05783_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_2 _11866_ (.A0(\core.cpuregs[28][14] ),
    .A1(_05367_),
    .S(_05779_),
    .X(_05784_));
 sky130_fd_sc_hd__buf_1 _11867_ (.A(_05784_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_2 _11868_ (.A0(\core.cpuregs[28][15] ),
    .A1(_05372_),
    .S(_05779_),
    .X(_05785_));
 sky130_fd_sc_hd__buf_1 _11869_ (.A(_05785_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_2 _11870_ (.A0(\core.cpuregs[28][16] ),
    .A1(_05377_),
    .S(_05779_),
    .X(_05786_));
 sky130_fd_sc_hd__buf_1 _11871_ (.A(_05786_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_2 _11872_ (.A0(\core.cpuregs[28][17] ),
    .A1(_05383_),
    .S(_05779_),
    .X(_05787_));
 sky130_fd_sc_hd__buf_1 _11873_ (.A(_05787_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_2 _11874_ (.A0(\core.cpuregs[28][18] ),
    .A1(_05388_),
    .S(_05779_),
    .X(_05788_));
 sky130_fd_sc_hd__buf_1 _11875_ (.A(_05788_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_2 _11876_ (.A0(\core.cpuregs[28][19] ),
    .A1(_05393_),
    .S(_05779_),
    .X(_05789_));
 sky130_fd_sc_hd__buf_1 _11877_ (.A(_05789_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_1 _11878_ (.A(_05767_),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_2 _11879_ (.A0(\core.cpuregs[28][20] ),
    .A1(_05399_),
    .S(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__buf_1 _11880_ (.A(_05791_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_2 _11881_ (.A0(\core.cpuregs[28][21] ),
    .A1(_05405_),
    .S(_05790_),
    .X(_05792_));
 sky130_fd_sc_hd__buf_1 _11882_ (.A(_05792_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_2 _11883_ (.A0(\core.cpuregs[28][22] ),
    .A1(_05410_),
    .S(_05790_),
    .X(_05793_));
 sky130_fd_sc_hd__buf_1 _11884_ (.A(_05793_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_2 _11885_ (.A0(\core.cpuregs[28][23] ),
    .A1(_05416_),
    .S(_05790_),
    .X(_05794_));
 sky130_fd_sc_hd__buf_1 _11886_ (.A(_05794_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_2 _11887_ (.A0(\core.cpuregs[28][24] ),
    .A1(_05421_),
    .S(_05790_),
    .X(_05795_));
 sky130_fd_sc_hd__buf_1 _11888_ (.A(_05795_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_2 _11889_ (.A0(\core.cpuregs[28][25] ),
    .A1(_05426_),
    .S(_05790_),
    .X(_05796_));
 sky130_fd_sc_hd__buf_1 _11890_ (.A(_05796_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_2 _11891_ (.A0(\core.cpuregs[28][26] ),
    .A1(_05432_),
    .S(_05790_),
    .X(_05797_));
 sky130_fd_sc_hd__buf_1 _11892_ (.A(_05797_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_2 _11893_ (.A0(\core.cpuregs[28][27] ),
    .A1(_05437_),
    .S(_05790_),
    .X(_05798_));
 sky130_fd_sc_hd__buf_1 _11894_ (.A(_05798_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_2 _11895_ (.A0(\core.cpuregs[28][28] ),
    .A1(_05442_),
    .S(_05790_),
    .X(_05799_));
 sky130_fd_sc_hd__buf_1 _11896_ (.A(_05799_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_2 _11897_ (.A0(\core.cpuregs[28][29] ),
    .A1(_05448_),
    .S(_05790_),
    .X(_05800_));
 sky130_fd_sc_hd__buf_1 _11898_ (.A(_05800_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_2 _11899_ (.A0(\core.cpuregs[28][30] ),
    .A1(_05453_),
    .S(_05767_),
    .X(_05801_));
 sky130_fd_sc_hd__buf_1 _11900_ (.A(_05801_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_2 _11901_ (.A0(\core.cpuregs[28][31] ),
    .A1(_05458_),
    .S(_05767_),
    .X(_05802_));
 sky130_fd_sc_hd__buf_1 _11902_ (.A(_05802_),
    .X(_00502_));
 sky130_fd_sc_hd__nand3_2 _11903_ (.A(\core.mem_do_rinst ),
    .B(_02024_),
    .C(_02029_),
    .Y(_05803_));
 sky130_fd_sc_hd__mux2_2 _11904_ (.A0(\core.mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(_02026_),
    .X(_05804_));
 sky130_fd_sc_hd__buf_1 _11905_ (.A(_05804_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_2 _11906_ (.A0(\core.mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(_03176_),
    .X(_05805_));
 sky130_fd_sc_hd__buf_1 _11907_ (.A(_05805_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_2 _11908_ (.A0(\core.mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(_02026_),
    .X(_05806_));
 sky130_fd_sc_hd__buf_1 _11909_ (.A(_05806_),
    .X(_01348_));
 sky130_fd_sc_hd__and3b_2 _11910_ (.A_N(_01349_),
    .B(_01347_),
    .C(_01348_),
    .X(_05807_));
 sky130_fd_sc_hd__mux2_2 _11911_ (.A0(\core.mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(_02026_),
    .X(_05808_));
 sky130_fd_sc_hd__buf_1 _11912_ (.A(_05808_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_2 _11913_ (.A0(\core.mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(_02026_),
    .X(_05809_));
 sky130_fd_sc_hd__buf_1 _11914_ (.A(_05809_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_2 _11915_ (.A0(\core.mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(_02026_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_1 _11916_ (.A(_05810_),
    .X(_01343_));
 sky130_fd_sc_hd__and3_2 _11917_ (.A(_02448_),
    .B(_01344_),
    .C(_01343_),
    .X(_05811_));
 sky130_fd_sc_hd__or2b_2 _11918_ (.A(_01346_),
    .B_N(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__mux2_2 _11919_ (.A0(\core.mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(_03176_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_1 _11920_ (.A(_05813_),
    .X(_01345_));
 sky130_fd_sc_hd__nor2_2 _11921_ (.A(_05812_),
    .B(_01345_),
    .Y(_05814_));
 sky130_fd_sc_hd__a22o_2 _11922_ (.A1(\core.is_alu_reg_reg ),
    .A2(_05803_),
    .B1(_05807_),
    .B2(_05814_),
    .X(_00503_));
 sky130_fd_sc_hd__nor3b_2 _11923_ (.A(_01349_),
    .B(_01348_),
    .C_N(_01347_),
    .Y(_05815_));
 sky130_fd_sc_hd__a22o_2 _11924_ (.A1(\core.is_alu_reg_imm ),
    .A2(_05803_),
    .B1(_05814_),
    .B2(_05815_),
    .X(_00504_));
 sky130_fd_sc_hd__and2b_2 _11925_ (.A_N(_05812_),
    .B(_01345_),
    .X(_05816_));
 sky130_fd_sc_hd__a22o_2 _11926_ (.A1(\core.instr_auipc ),
    .A2(_05803_),
    .B1(_05815_),
    .B2(_05816_),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_2 _11927_ (.A1(\core.instr_lui ),
    .A2(_05803_),
    .B1(_05807_),
    .B2(_05816_),
    .X(_00506_));
 sky130_fd_sc_hd__o21ai_2 _11928_ (.A1(\core.cpu_state[1] ),
    .A2(_02045_),
    .B1(_02046_),
    .Y(_05817_));
 sky130_fd_sc_hd__a22o_2 _11929_ (.A1(\core.instr_lb ),
    .A2(_02051_),
    .B1(_05817_),
    .B2(\core.latched_is_lb ),
    .X(_05818_));
 sky130_fd_sc_hd__and2_2 _11930_ (.A(_04144_),
    .B(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__buf_1 _11931_ (.A(_05819_),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_2 _11932_ (.A1(\core.instr_lh ),
    .A2(_02051_),
    .B1(_05817_),
    .B2(\core.latched_is_lh ),
    .X(_05820_));
 sky130_fd_sc_hd__and2_2 _11933_ (.A(_04144_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_1 _11934_ (.A(_05821_),
    .X(_00508_));
 sky130_fd_sc_hd__o21a_2 _11935_ (.A1(_02117_),
    .A2(_02445_),
    .B1(_02450_),
    .X(_05822_));
 sky130_fd_sc_hd__o21ai_2 _11936_ (.A1(_02236_),
    .A2(\core.instr_jalr ),
    .B1(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__nor2_2 _11937_ (.A(\core.latched_branch ),
    .B(_02079_),
    .Y(_05824_));
 sky130_fd_sc_hd__a211o_2 _11938_ (.A1(_02079_),
    .A2(_03672_),
    .B1(_05824_),
    .C1(_02450_),
    .X(_05825_));
 sky130_fd_sc_hd__a21oi_2 _11939_ (.A1(_05823_),
    .A2(_05825_),
    .B1(_02055_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_2 _11940_ (.A(_02234_),
    .B(_02079_),
    .Y(_05826_));
 sky130_fd_sc_hd__o2bb2a_2 _11941_ (.A1_N(_03862_),
    .A2_N(_05826_),
    .B1(_02236_),
    .B2(_02234_),
    .X(_05827_));
 sky130_fd_sc_hd__nor2_2 _11942_ (.A(_02055_),
    .B(_05827_),
    .Y(_00511_));
 sky130_fd_sc_hd__nor2_2 _11943_ (.A(_02055_),
    .B(_02076_),
    .Y(_00512_));
 sky130_fd_sc_hd__or2_2 _11944_ (.A(_02108_),
    .B(\core.decoder_pseudo_trigger ),
    .X(_05828_));
 sky130_fd_sc_hd__buf_1 _11945_ (.A(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__buf_1 _11946_ (.A(_05828_),
    .X(_05830_));
 sky130_fd_sc_hd__or2b_2 _11947_ (.A(\core.mem_rdata_q[13] ),
    .B_N(\core.mem_rdata_q[12] ),
    .X(_05831_));
 sky130_fd_sc_hd__or2_2 _11948_ (.A(\core.mem_rdata_q[14] ),
    .B(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__nor2_2 _11949_ (.A(_05830_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__a22o_2 _11950_ (.A1(\core.instr_bne ),
    .A2(_05829_),
    .B1(_05833_),
    .B2(_02236_),
    .X(_05834_));
 sky130_fd_sc_hd__and2_2 _11951_ (.A(_04144_),
    .B(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__buf_1 _11952_ (.A(_05835_),
    .X(_00513_));
 sky130_fd_sc_hd__or3b_2 _11953_ (.A(_05462_),
    .B(\core.latched_rd[1] ),
    .C_N(\core.latched_rd[0] ),
    .X(_05836_));
 sky130_fd_sc_hd__buf_1 _11954_ (.A(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__nor2_2 _11955_ (.A(_05285_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__buf_1 _11956_ (.A(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_2 _11957_ (.A0(\core.cpuregs[21][0] ),
    .A1(_05284_),
    .S(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__buf_1 _11958_ (.A(_05840_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_2 _11959_ (.A0(\core.cpuregs[21][1] ),
    .A1(_05292_),
    .S(_05839_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_1 _11960_ (.A(_05841_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_2 _11961_ (.A0(\core.cpuregs[21][2] ),
    .A1(_05297_),
    .S(_05839_),
    .X(_05842_));
 sky130_fd_sc_hd__buf_1 _11962_ (.A(_05842_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_2 _11963_ (.A0(\core.cpuregs[21][3] ),
    .A1(_05304_),
    .S(_05839_),
    .X(_05843_));
 sky130_fd_sc_hd__buf_1 _11964_ (.A(_05843_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_2 _11965_ (.A0(\core.cpuregs[21][4] ),
    .A1(_05310_),
    .S(_05839_),
    .X(_05844_));
 sky130_fd_sc_hd__buf_1 _11966_ (.A(_05844_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_2 _11967_ (.A0(\core.cpuregs[21][5] ),
    .A1(_05315_),
    .S(_05839_),
    .X(_05845_));
 sky130_fd_sc_hd__buf_1 _11968_ (.A(_05845_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_2 _11969_ (.A0(\core.cpuregs[21][6] ),
    .A1(_05320_),
    .S(_05839_),
    .X(_05846_));
 sky130_fd_sc_hd__buf_1 _11970_ (.A(_05846_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_2 _11971_ (.A0(\core.cpuregs[21][7] ),
    .A1(_05326_),
    .S(_05839_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _11972_ (.A(_05847_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_2 _11973_ (.A0(\core.cpuregs[21][8] ),
    .A1(_05332_),
    .S(_05839_),
    .X(_05848_));
 sky130_fd_sc_hd__buf_1 _11974_ (.A(_05848_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_2 _11975_ (.A0(\core.cpuregs[21][9] ),
    .A1(_05337_),
    .S(_05839_),
    .X(_05849_));
 sky130_fd_sc_hd__buf_1 _11976_ (.A(_05849_),
    .X(_00523_));
 sky130_fd_sc_hd__buf_1 _11977_ (.A(_05838_),
    .X(_05850_));
 sky130_fd_sc_hd__mux2_2 _11978_ (.A0(\core.cpuregs[21][10] ),
    .A1(_05343_),
    .S(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__buf_1 _11979_ (.A(_05851_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_2 _11980_ (.A0(\core.cpuregs[21][11] ),
    .A1(_05349_),
    .S(_05850_),
    .X(_05852_));
 sky130_fd_sc_hd__buf_1 _11981_ (.A(_05852_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_2 _11982_ (.A0(\core.cpuregs[21][12] ),
    .A1(_05355_),
    .S(_05850_),
    .X(_05853_));
 sky130_fd_sc_hd__buf_1 _11983_ (.A(_05853_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_2 _11984_ (.A0(\core.cpuregs[21][13] ),
    .A1(_05360_),
    .S(_05850_),
    .X(_05854_));
 sky130_fd_sc_hd__buf_1 _11985_ (.A(_05854_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_2 _11986_ (.A0(\core.cpuregs[21][14] ),
    .A1(_05367_),
    .S(_05850_),
    .X(_05855_));
 sky130_fd_sc_hd__buf_1 _11987_ (.A(_05855_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_2 _11988_ (.A0(\core.cpuregs[21][15] ),
    .A1(_05372_),
    .S(_05850_),
    .X(_05856_));
 sky130_fd_sc_hd__buf_1 _11989_ (.A(_05856_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_2 _11990_ (.A0(\core.cpuregs[21][16] ),
    .A1(_05377_),
    .S(_05850_),
    .X(_05857_));
 sky130_fd_sc_hd__buf_1 _11991_ (.A(_05857_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_2 _11992_ (.A0(\core.cpuregs[21][17] ),
    .A1(_05383_),
    .S(_05850_),
    .X(_05858_));
 sky130_fd_sc_hd__buf_1 _11993_ (.A(_05858_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_2 _11994_ (.A0(\core.cpuregs[21][18] ),
    .A1(_05388_),
    .S(_05850_),
    .X(_05859_));
 sky130_fd_sc_hd__buf_1 _11995_ (.A(_05859_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_2 _11996_ (.A0(\core.cpuregs[21][19] ),
    .A1(_05393_),
    .S(_05850_),
    .X(_05860_));
 sky130_fd_sc_hd__buf_1 _11997_ (.A(_05860_),
    .X(_00533_));
 sky130_fd_sc_hd__buf_1 _11998_ (.A(_05838_),
    .X(_05861_));
 sky130_fd_sc_hd__mux2_2 _11999_ (.A0(\core.cpuregs[21][20] ),
    .A1(_05399_),
    .S(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__buf_1 _12000_ (.A(_05862_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_2 _12001_ (.A0(\core.cpuregs[21][21] ),
    .A1(_05405_),
    .S(_05861_),
    .X(_05863_));
 sky130_fd_sc_hd__buf_1 _12002_ (.A(_05863_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_2 _12003_ (.A0(\core.cpuregs[21][22] ),
    .A1(_05410_),
    .S(_05861_),
    .X(_05864_));
 sky130_fd_sc_hd__buf_1 _12004_ (.A(_05864_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_2 _12005_ (.A0(\core.cpuregs[21][23] ),
    .A1(_05416_),
    .S(_05861_),
    .X(_05865_));
 sky130_fd_sc_hd__buf_1 _12006_ (.A(_05865_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_2 _12007_ (.A0(\core.cpuregs[21][24] ),
    .A1(_05421_),
    .S(_05861_),
    .X(_05866_));
 sky130_fd_sc_hd__buf_1 _12008_ (.A(_05866_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_2 _12009_ (.A0(\core.cpuregs[21][25] ),
    .A1(_05426_),
    .S(_05861_),
    .X(_05867_));
 sky130_fd_sc_hd__buf_1 _12010_ (.A(_05867_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_2 _12011_ (.A0(\core.cpuregs[21][26] ),
    .A1(_05432_),
    .S(_05861_),
    .X(_05868_));
 sky130_fd_sc_hd__buf_1 _12012_ (.A(_05868_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_2 _12013_ (.A0(\core.cpuregs[21][27] ),
    .A1(_05437_),
    .S(_05861_),
    .X(_05869_));
 sky130_fd_sc_hd__buf_1 _12014_ (.A(_05869_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_2 _12015_ (.A0(\core.cpuregs[21][28] ),
    .A1(_05442_),
    .S(_05861_),
    .X(_05870_));
 sky130_fd_sc_hd__buf_1 _12016_ (.A(_05870_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_2 _12017_ (.A0(\core.cpuregs[21][29] ),
    .A1(_05448_),
    .S(_05861_),
    .X(_05871_));
 sky130_fd_sc_hd__buf_1 _12018_ (.A(_05871_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_2 _12019_ (.A0(\core.cpuregs[21][30] ),
    .A1(_05453_),
    .S(_05838_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _12020_ (.A(_05872_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_2 _12021_ (.A0(\core.cpuregs[21][31] ),
    .A1(_05458_),
    .S(_05838_),
    .X(_05873_));
 sky130_fd_sc_hd__buf_1 _12022_ (.A(_05873_),
    .X(_00545_));
 sky130_fd_sc_hd__and3b_2 _12023_ (.A_N(_01347_),
    .B(_01348_),
    .C(_01349_),
    .X(_05874_));
 sky130_fd_sc_hd__and3_2 _12024_ (.A(_01346_),
    .B(_01345_),
    .C(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__a22o_2 _12025_ (.A1(_02019_),
    .A2(_05803_),
    .B1(_05811_),
    .B2(_05875_),
    .X(_00546_));
 sky130_fd_sc_hd__nor2_2 _12026_ (.A(_02108_),
    .B(\core.decoder_pseudo_trigger ),
    .Y(_05876_));
 sky130_fd_sc_hd__buf_1 _12027_ (.A(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__inv_2 _12028_ (.A(\core.mem_rdata_q[14] ),
    .Y(_05878_));
 sky130_fd_sc_hd__nor2_2 _12029_ (.A(\core.mem_rdata_q[12] ),
    .B(\core.mem_rdata_q[13] ),
    .Y(_05879_));
 sky130_fd_sc_hd__and2_2 _12030_ (.A(_05878_),
    .B(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__and2_2 _12031_ (.A(_05877_),
    .B(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__a22o_2 _12032_ (.A1(\core.instr_beq ),
    .A2(_05829_),
    .B1(_05881_),
    .B2(_02236_),
    .X(_05882_));
 sky130_fd_sc_hd__and2_2 _12033_ (.A(_04144_),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__buf_1 _12034_ (.A(_05883_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_2 _12035_ (.A(_05464_),
    .B(_05657_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _12036_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__mux2_2 _12037_ (.A0(_05460_),
    .A1(\core.cpuregs[26][0] ),
    .S(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__buf_1 _12038_ (.A(_05886_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_2 _12039_ (.A0(_05468_),
    .A1(\core.cpuregs[26][1] ),
    .S(_05885_),
    .X(_05887_));
 sky130_fd_sc_hd__buf_1 _12040_ (.A(_05887_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_2 _12041_ (.A0(_05470_),
    .A1(\core.cpuregs[26][2] ),
    .S(_05885_),
    .X(_05888_));
 sky130_fd_sc_hd__buf_1 _12042_ (.A(_05888_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_2 _12043_ (.A0(_05472_),
    .A1(\core.cpuregs[26][3] ),
    .S(_05885_),
    .X(_05889_));
 sky130_fd_sc_hd__buf_1 _12044_ (.A(_05889_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_2 _12045_ (.A0(_05474_),
    .A1(\core.cpuregs[26][4] ),
    .S(_05885_),
    .X(_05890_));
 sky130_fd_sc_hd__buf_1 _12046_ (.A(_05890_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_2 _12047_ (.A0(_05476_),
    .A1(\core.cpuregs[26][5] ),
    .S(_05885_),
    .X(_05891_));
 sky130_fd_sc_hd__buf_1 _12048_ (.A(_05891_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_2 _12049_ (.A0(_05478_),
    .A1(\core.cpuregs[26][6] ),
    .S(_05885_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _12050_ (.A(_05892_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_2 _12051_ (.A0(_05480_),
    .A1(\core.cpuregs[26][7] ),
    .S(_05885_),
    .X(_05893_));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_05893_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_2 _12053_ (.A0(_05482_),
    .A1(\core.cpuregs[26][8] ),
    .S(_05885_),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _12054_ (.A(_05894_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_2 _12055_ (.A0(_05484_),
    .A1(\core.cpuregs[26][9] ),
    .S(_05885_),
    .X(_05895_));
 sky130_fd_sc_hd__buf_1 _12056_ (.A(_05895_),
    .X(_00557_));
 sky130_fd_sc_hd__buf_1 _12057_ (.A(_05884_),
    .X(_05896_));
 sky130_fd_sc_hd__mux2_2 _12058_ (.A0(_05486_),
    .A1(\core.cpuregs[26][10] ),
    .S(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__buf_1 _12059_ (.A(_05897_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_2 _12060_ (.A0(_05489_),
    .A1(\core.cpuregs[26][11] ),
    .S(_05896_),
    .X(_05898_));
 sky130_fd_sc_hd__buf_1 _12061_ (.A(_05898_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_2 _12062_ (.A0(_05491_),
    .A1(\core.cpuregs[26][12] ),
    .S(_05896_),
    .X(_05899_));
 sky130_fd_sc_hd__buf_1 _12063_ (.A(_05899_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_2 _12064_ (.A0(_05493_),
    .A1(\core.cpuregs[26][13] ),
    .S(_05896_),
    .X(_05900_));
 sky130_fd_sc_hd__buf_1 _12065_ (.A(_05900_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_2 _12066_ (.A0(_05495_),
    .A1(\core.cpuregs[26][14] ),
    .S(_05896_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_1 _12067_ (.A(_05901_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_2 _12068_ (.A0(_05497_),
    .A1(\core.cpuregs[26][15] ),
    .S(_05896_),
    .X(_05902_));
 sky130_fd_sc_hd__buf_1 _12069_ (.A(_05902_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_2 _12070_ (.A0(_05499_),
    .A1(\core.cpuregs[26][16] ),
    .S(_05896_),
    .X(_05903_));
 sky130_fd_sc_hd__buf_1 _12071_ (.A(_05903_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_2 _12072_ (.A0(_05501_),
    .A1(\core.cpuregs[26][17] ),
    .S(_05896_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_1 _12073_ (.A(_05904_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_2 _12074_ (.A0(_05503_),
    .A1(\core.cpuregs[26][18] ),
    .S(_05896_),
    .X(_05905_));
 sky130_fd_sc_hd__buf_1 _12075_ (.A(_05905_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_2 _12076_ (.A0(_05505_),
    .A1(\core.cpuregs[26][19] ),
    .S(_05896_),
    .X(_05906_));
 sky130_fd_sc_hd__buf_1 _12077_ (.A(_05906_),
    .X(_00567_));
 sky130_fd_sc_hd__buf_1 _12078_ (.A(_05884_),
    .X(_05907_));
 sky130_fd_sc_hd__mux2_2 _12079_ (.A0(_05507_),
    .A1(\core.cpuregs[26][20] ),
    .S(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__buf_1 _12080_ (.A(_05908_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_2 _12081_ (.A0(_05510_),
    .A1(\core.cpuregs[26][21] ),
    .S(_05907_),
    .X(_05909_));
 sky130_fd_sc_hd__buf_1 _12082_ (.A(_05909_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_2 _12083_ (.A0(_05512_),
    .A1(\core.cpuregs[26][22] ),
    .S(_05907_),
    .X(_05910_));
 sky130_fd_sc_hd__buf_1 _12084_ (.A(_05910_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_2 _12085_ (.A0(_05514_),
    .A1(\core.cpuregs[26][23] ),
    .S(_05907_),
    .X(_05911_));
 sky130_fd_sc_hd__buf_1 _12086_ (.A(_05911_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_2 _12087_ (.A0(_05516_),
    .A1(\core.cpuregs[26][24] ),
    .S(_05907_),
    .X(_05912_));
 sky130_fd_sc_hd__buf_1 _12088_ (.A(_05912_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_2 _12089_ (.A0(_05518_),
    .A1(\core.cpuregs[26][25] ),
    .S(_05907_),
    .X(_05913_));
 sky130_fd_sc_hd__buf_1 _12090_ (.A(_05913_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_2 _12091_ (.A0(_05520_),
    .A1(\core.cpuregs[26][26] ),
    .S(_05907_),
    .X(_05914_));
 sky130_fd_sc_hd__buf_1 _12092_ (.A(_05914_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_2 _12093_ (.A0(_05522_),
    .A1(\core.cpuregs[26][27] ),
    .S(_05907_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_1 _12094_ (.A(_05915_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_2 _12095_ (.A0(_05524_),
    .A1(\core.cpuregs[26][28] ),
    .S(_05907_),
    .X(_05916_));
 sky130_fd_sc_hd__buf_1 _12096_ (.A(_05916_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_2 _12097_ (.A0(_05526_),
    .A1(\core.cpuregs[26][29] ),
    .S(_05907_),
    .X(_05917_));
 sky130_fd_sc_hd__buf_1 _12098_ (.A(_05917_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_2 _12099_ (.A0(_05528_),
    .A1(\core.cpuregs[26][30] ),
    .S(_05884_),
    .X(_05918_));
 sky130_fd_sc_hd__buf_1 _12100_ (.A(_05918_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_2 _12101_ (.A0(_05530_),
    .A1(\core.cpuregs[26][31] ),
    .S(_05884_),
    .X(_05919_));
 sky130_fd_sc_hd__buf_1 _12102_ (.A(_05919_),
    .X(_00579_));
 sky130_fd_sc_hd__buf_1 _12103_ (.A(_05830_),
    .X(_05920_));
 sky130_fd_sc_hd__buf_1 _12104_ (.A(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__a22o_2 _12105_ (.A1(\core.instr_sh ),
    .A2(_05921_),
    .B1(_05833_),
    .B2(_02090_),
    .X(_00580_));
 sky130_fd_sc_hd__or3b_2 _12106_ (.A(\core.mem_rdata_q[12] ),
    .B(\core.mem_rdata_q[14] ),
    .C_N(\core.mem_rdata_q[13] ),
    .X(_05922_));
 sky130_fd_sc_hd__inv_2 _12107_ (.A(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__and2_2 _12108_ (.A(\core.is_alu_reg_imm ),
    .B(_05876_),
    .X(_05924_));
 sky130_fd_sc_hd__buf_1 _12109_ (.A(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a22o_2 _12110_ (.A1(\core.instr_slti ),
    .A2(_05829_),
    .B1(_05923_),
    .B2(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__and2_2 _12111_ (.A(_04144_),
    .B(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__buf_1 _12112_ (.A(_05927_),
    .X(_00581_));
 sky130_fd_sc_hd__buf_1 _12113_ (.A(_02052_),
    .X(_05928_));
 sky130_fd_sc_hd__and3_2 _12114_ (.A(\core.mem_rdata_q[12] ),
    .B(\core.mem_rdata_q[13] ),
    .C(_05878_),
    .X(_05929_));
 sky130_fd_sc_hd__a22o_2 _12115_ (.A1(\core.instr_sltiu ),
    .A2(_05829_),
    .B1(_05925_),
    .B2(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__and2_2 _12116_ (.A(_05928_),
    .B(_05930_),
    .X(_05931_));
 sky130_fd_sc_hd__buf_1 _12117_ (.A(_05931_),
    .X(_00582_));
 sky130_fd_sc_hd__buf_1 _12118_ (.A(_05828_),
    .X(_05932_));
 sky130_fd_sc_hd__and3b_2 _12119_ (.A_N(\core.mem_rdata_q[12] ),
    .B(\core.mem_rdata_q[13] ),
    .C(\core.mem_rdata_q[14] ),
    .X(_05933_));
 sky130_fd_sc_hd__a22o_2 _12120_ (.A1(\core.instr_ori ),
    .A2(_05932_),
    .B1(_05925_),
    .B2(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__and2_2 _12121_ (.A(_05928_),
    .B(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__buf_1 _12122_ (.A(_05935_),
    .X(_00583_));
 sky130_fd_sc_hd__or2_2 _12123_ (.A(\core.cpu_state[1] ),
    .B(_02488_),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_2 _12124_ (.A0(_02057_),
    .A1(_05936_),
    .S(_02056_),
    .X(_05937_));
 sky130_fd_sc_hd__or4b_2 _12125_ (.A(\core.cpu_state[2] ),
    .B(_02116_),
    .C(_02087_),
    .D_N(_05936_),
    .X(_05938_));
 sky130_fd_sc_hd__o221a_2 _12126_ (.A1(\core.latched_store ),
    .A2(_05937_),
    .B1(_05938_),
    .B2(_05822_),
    .C1(_03680_),
    .X(_00584_));
 sky130_fd_sc_hd__or3_2 _12127_ (.A(\core.mem_rdata_q[25] ),
    .B(\core.mem_rdata_q[26] ),
    .C(\core.mem_rdata_q[27] ),
    .X(_05939_));
 sky130_fd_sc_hd__nor4_2 _12128_ (.A(\core.mem_rdata_q[28] ),
    .B(\core.mem_rdata_q[29] ),
    .C(\core.mem_rdata_q[31] ),
    .D(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__or2b_2 _12129_ (.A(\core.mem_rdata_q[30] ),
    .B_N(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__nor2_2 _12130_ (.A(_05831_),
    .B(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__buf_1 _12131_ (.A(_05829_),
    .X(_05943_));
 sky130_fd_sc_hd__a32o_2 _12132_ (.A1(\core.mem_rdata_q[14] ),
    .A2(_05925_),
    .A3(_05942_),
    .B1(_05943_),
    .B2(\core.instr_srli ),
    .X(_00585_));
 sky130_fd_sc_hd__nand2_2 _12133_ (.A(\core.is_alu_reg_reg ),
    .B(_05877_),
    .Y(_05944_));
 sky130_fd_sc_hd__nor2_2 _12134_ (.A(_05941_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__a22o_2 _12135_ (.A1(\core.instr_add ),
    .A2(_05932_),
    .B1(_05880_),
    .B2(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__and2_2 _12136_ (.A(_05928_),
    .B(_05946_),
    .X(_05947_));
 sky130_fd_sc_hd__buf_1 _12137_ (.A(_05947_),
    .X(_00586_));
 sky130_fd_sc_hd__or2_2 _12138_ (.A(_05941_),
    .B(_05944_),
    .X(_05948_));
 sky130_fd_sc_hd__o2bb2a_2 _12139_ (.A1_N(\core.instr_sll ),
    .A2_N(_05920_),
    .B1(_05832_),
    .B2(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__nor2_2 _12140_ (.A(_02055_),
    .B(_05949_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_2 _12141_ (.A(\core.mem_rdata_q[14] ),
    .B(_05879_),
    .Y(_05950_));
 sky130_fd_sc_hd__o2bb2a_2 _12142_ (.A1_N(\core.instr_xor ),
    .A2_N(_05920_),
    .B1(_05948_),
    .B2(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__nor2_2 _12143_ (.A(_02055_),
    .B(_05951_),
    .Y(_00588_));
 sky130_fd_sc_hd__and2_2 _12144_ (.A(\core.is_alu_reg_reg ),
    .B(_05876_),
    .X(_05952_));
 sky130_fd_sc_hd__nor2_2 _12145_ (.A(_05878_),
    .B(_05831_),
    .Y(_05953_));
 sky130_fd_sc_hd__and3_2 _12146_ (.A(\core.mem_rdata_q[30] ),
    .B(_05940_),
    .C(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__a22o_2 _12147_ (.A1(\core.instr_sra ),
    .A2(_05932_),
    .B1(_05952_),
    .B2(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__and2_2 _12148_ (.A(_05928_),
    .B(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_1 _12149_ (.A(_05956_),
    .X(_00589_));
 sky130_fd_sc_hd__or4_2 _12150_ (.A(\core.instr_slt ),
    .B(\core.instr_sltu ),
    .C(_02236_),
    .D(\core.instr_slti ),
    .X(_05957_));
 sky130_fd_sc_hd__o211a_2 _12151_ (.A1(\core.instr_sltiu ),
    .A2(_05957_),
    .B1(_05921_),
    .C1(_03665_),
    .X(_00590_));
 sky130_fd_sc_hd__nand2_2 _12152_ (.A(_02236_),
    .B(_02450_),
    .Y(_05958_));
 sky130_fd_sc_hd__a21o_2 _12153_ (.A1(_05958_),
    .A2(_05826_),
    .B1(_02049_),
    .X(_05959_));
 sky130_fd_sc_hd__nor2_2 _12154_ (.A(_02523_),
    .B(_03791_),
    .Y(_05960_));
 sky130_fd_sc_hd__a22o_2 _12155_ (.A1(\core.latched_rd[0] ),
    .A2(_05959_),
    .B1(_05960_),
    .B2(\core.decoded_rd[0] ),
    .X(_00591_));
 sky130_fd_sc_hd__a22o_2 _12156_ (.A1(\core.latched_rd[1] ),
    .A2(_05959_),
    .B1(_05960_),
    .B2(\core.decoded_rd[1] ),
    .X(_00592_));
 sky130_fd_sc_hd__a22o_2 _12157_ (.A1(\core.latched_rd[2] ),
    .A2(_05959_),
    .B1(_05960_),
    .B2(\core.decoded_rd[2] ),
    .X(_00593_));
 sky130_fd_sc_hd__a22o_2 _12158_ (.A1(\core.latched_rd[3] ),
    .A2(_05959_),
    .B1(_05960_),
    .B2(\core.decoded_rd[3] ),
    .X(_00594_));
 sky130_fd_sc_hd__a22o_2 _12159_ (.A1(\core.latched_rd[4] ),
    .A2(_05959_),
    .B1(_05960_),
    .B2(\core.decoded_rd[4] ),
    .X(_00595_));
 sky130_fd_sc_hd__o21a_2 _12160_ (.A1(_02466_),
    .A2(_03212_),
    .B1(_03210_),
    .X(_05961_));
 sky130_fd_sc_hd__o22a_2 _12161_ (.A1(mem_wstrb[0]),
    .A2(_03214_),
    .B1(_05269_),
    .B2(_05961_),
    .X(_00596_));
 sky130_fd_sc_hd__and2b_2 _12162_ (.A_N(_05269_),
    .B(_03210_),
    .X(_05962_));
 sky130_fd_sc_hd__nor2_2 _12163_ (.A(_02123_),
    .B(_02070_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_2 _12164_ (.A1(_02476_),
    .A2(_05963_),
    .B1(_02472_),
    .Y(_05964_));
 sky130_fd_sc_hd__mux2_2 _12165_ (.A0(_05964_),
    .A1(mem_wstrb[1]),
    .S(_03212_),
    .X(_05965_));
 sky130_fd_sc_hd__a22o_2 _12166_ (.A1(mem_wstrb[1]),
    .A2(_05269_),
    .B1(_05962_),
    .B2(_05965_),
    .X(_00597_));
 sky130_fd_sc_hd__o31a_2 _12167_ (.A1(_05704_),
    .A2(_02469_),
    .A3(_03212_),
    .B1(_03210_),
    .X(_05966_));
 sky130_fd_sc_hd__o22a_2 _12168_ (.A1(mem_wstrb[2]),
    .A2(_03214_),
    .B1(_05269_),
    .B2(_05966_),
    .X(_00598_));
 sky130_fd_sc_hd__o21ai_2 _12169_ (.A1(_02365_),
    .A2(_05963_),
    .B1(_02472_),
    .Y(_05967_));
 sky130_fd_sc_hd__mux2_2 _12170_ (.A0(_05967_),
    .A1(mem_wstrb[3]),
    .S(_03212_),
    .X(_05968_));
 sky130_fd_sc_hd__a22o_2 _12171_ (.A1(mem_wstrb[3]),
    .A2(_05269_),
    .B1(_05962_),
    .B2(_05968_),
    .X(_00599_));
 sky130_fd_sc_hd__nor4b_2 _12172_ (.A(\core.mem_rdata_q[24] ),
    .B(\core.mem_rdata_q[25] ),
    .C(\core.mem_rdata_q[26] ),
    .D_N(\core.mem_rdata_q[27] ),
    .Y(_05969_));
 sky130_fd_sc_hd__or3_2 _12173_ (.A(\core.mem_rdata_q[22] ),
    .B(\core.mem_rdata_q[23] ),
    .C(_05830_),
    .X(_05970_));
 sky130_fd_sc_hd__nor2_2 _12174_ (.A(\core.mem_rdata_q[21] ),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__and4b_2 _12175_ (.A_N(\core.mem_rdata_q[3] ),
    .B(\core.mem_rdata_q[4] ),
    .C(\core.mem_rdata_q[5] ),
    .D(\core.mem_rdata_q[6] ),
    .X(_05972_));
 sky130_fd_sc_hd__nor4_2 _12176_ (.A(\core.mem_rdata_q[17] ),
    .B(\core.mem_rdata_q[18] ),
    .C(\core.mem_rdata_q[19] ),
    .D(\core.mem_rdata_q[2] ),
    .Y(_05973_));
 sky130_fd_sc_hd__nor3_2 _12177_ (.A(\core.mem_rdata_q[28] ),
    .B(\core.mem_rdata_q[15] ),
    .C(\core.mem_rdata_q[16] ),
    .Y(_05974_));
 sky130_fd_sc_hd__and4b_2 _12178_ (.A_N(\core.mem_rdata_q[29] ),
    .B(\core.mem_rdata_q[30] ),
    .C(\core.mem_rdata_q[0] ),
    .D(\core.mem_rdata_q[1] ),
    .X(_05975_));
 sky130_fd_sc_hd__and3_2 _12179_ (.A(\core.mem_rdata_q[31] ),
    .B(_05974_),
    .C(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__and4_2 _12180_ (.A(_05923_),
    .B(_05972_),
    .C(_05973_),
    .D(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__a32o_2 _12181_ (.A1(_05969_),
    .A2(_05971_),
    .A3(_05977_),
    .B1(_05943_),
    .B2(_02532_),
    .X(_00600_));
 sky130_fd_sc_hd__o221ai_2 _12182_ (.A1(_05271_),
    .A2(_05269_),
    .B1(_05274_),
    .B2(mem_ready),
    .C1(_05273_),
    .Y(_05978_));
 sky130_fd_sc_hd__a21o_2 _12183_ (.A1(mem_valid),
    .A2(_05978_),
    .B1(_03214_),
    .X(_00601_));
 sky130_fd_sc_hd__nor3_2 _12184_ (.A(\core.mem_rdata_q[4] ),
    .B(\core.mem_rdata_q[5] ),
    .C(\core.mem_rdata_q[6] ),
    .Y(_05979_));
 sky130_fd_sc_hd__and4_2 _12185_ (.A(\core.mem_rdata_q[0] ),
    .B(\core.mem_rdata_q[1] ),
    .C(\core.mem_rdata_q[2] ),
    .D(\core.mem_rdata_q[3] ),
    .X(_05980_));
 sky130_fd_sc_hd__a32o_2 _12186_ (.A1(_05881_),
    .A2(_05979_),
    .A3(_05980_),
    .B1(_05829_),
    .B2(\core.instr_fence ),
    .X(_05981_));
 sky130_fd_sc_hd__and2_2 _12187_ (.A(_05928_),
    .B(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__buf_1 _12188_ (.A(_05982_),
    .X(_00602_));
 sky130_fd_sc_hd__and3_2 _12189_ (.A(_02056_),
    .B(_02076_),
    .C(_03728_),
    .X(_05983_));
 sky130_fd_sc_hd__nor2_2 _12190_ (.A(_02048_),
    .B(_02029_),
    .Y(_05984_));
 sky130_fd_sc_hd__a32o_2 _12191_ (.A1(_02032_),
    .A2(_02454_),
    .A3(_05983_),
    .B1(_05984_),
    .B2(\core.mem_do_wdata ),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_2 _12192_ (.A0(\core.decoded_imm[0] ),
    .A1(_05554_),
    .S(_02095_),
    .X(_05985_));
 sky130_fd_sc_hd__nor2_2 _12193_ (.A(_02048_),
    .B(_02056_),
    .Y(_05986_));
 sky130_fd_sc_hd__buf_1 _12194_ (.A(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__mux2_2 _12195_ (.A0(_02368_),
    .A1(_05985_),
    .S(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__buf_1 _12196_ (.A(_05988_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_2 _12197_ (.A0(\core.decoded_imm[1] ),
    .A1(_05581_),
    .S(_02095_),
    .X(_05989_));
 sky130_fd_sc_hd__mux2_2 _12198_ (.A0(_02366_),
    .A1(_05989_),
    .S(_05987_),
    .X(_05990_));
 sky130_fd_sc_hd__buf_1 _12199_ (.A(_05990_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_2 _12200_ (.A0(\core.decoded_imm[2] ),
    .A1(_02176_),
    .S(_02095_),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_2 _12201_ (.A0(\core.mem_la_wdata[2] ),
    .A1(_05991_),
    .S(_05986_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_1 _12202_ (.A(_05992_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_2 _12203_ (.A0(\core.decoded_imm[3] ),
    .A1(_02206_),
    .S(_02095_),
    .X(_05993_));
 sky130_fd_sc_hd__mux2_2 _12204_ (.A0(\core.mem_la_wdata[3] ),
    .A1(_05993_),
    .S(_05986_),
    .X(_05994_));
 sky130_fd_sc_hd__buf_1 _12205_ (.A(_05994_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_2 _12206_ (.A0(\core.decoded_imm[4] ),
    .A1(_02232_),
    .S(_02095_),
    .X(_05995_));
 sky130_fd_sc_hd__mux2_2 _12207_ (.A0(\core.mem_la_wdata[4] ),
    .A1(_05995_),
    .S(_05986_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_1 _12208_ (.A(_05996_),
    .X(_00608_));
 sky130_fd_sc_hd__and2_2 _12209_ (.A(_02095_),
    .B(_02175_),
    .X(_05997_));
 sky130_fd_sc_hd__buf_1 _12210_ (.A(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__buf_1 _12211_ (.A(_02132_),
    .X(_05999_));
 sky130_fd_sc_hd__buf_1 _12212_ (.A(_02134_),
    .X(_06000_));
 sky130_fd_sc_hd__mux4_2 _12213_ (.A0(\core.cpuregs[12][5] ),
    .A1(\core.cpuregs[13][5] ),
    .A2(\core.cpuregs[14][5] ),
    .A3(\core.cpuregs[15][5] ),
    .S0(_06000_),
    .S1(_02159_),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_2 _12214_ (.A0(\core.cpuregs[8][5] ),
    .A1(\core.cpuregs[9][5] ),
    .S(_02149_),
    .X(_06002_));
 sky130_fd_sc_hd__mux2_2 _12215_ (.A0(\core.cpuregs[10][5] ),
    .A1(\core.cpuregs[11][5] ),
    .S(_02155_),
    .X(_06003_));
 sky130_fd_sc_hd__a21o_2 _12216_ (.A1(_02159_),
    .A2(_06003_),
    .B1(_02138_),
    .X(_06004_));
 sky130_fd_sc_hd__a21o_2 _12217_ (.A1(_02167_),
    .A2(_06002_),
    .B1(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__o211a_2 _12218_ (.A1(_05999_),
    .A2(_06001_),
    .B1(_06005_),
    .C1(_02152_),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_2 _12219_ (.A0(\core.cpuregs[4][5] ),
    .A1(\core.cpuregs[5][5] ),
    .S(_02149_),
    .X(_06007_));
 sky130_fd_sc_hd__and2_2 _12220_ (.A(_02167_),
    .B(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__mux2_2 _12221_ (.A0(\core.cpuregs[6][5] ),
    .A1(\core.cpuregs[7][5] ),
    .S(_02149_),
    .X(_06009_));
 sky130_fd_sc_hd__and2_2 _12222_ (.A(_02159_),
    .B(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__mux4_2 _12223_ (.A0(\core.cpuregs[0][5] ),
    .A1(\core.cpuregs[1][5] ),
    .A2(\core.cpuregs[2][5] ),
    .A3(\core.cpuregs[3][5] ),
    .S0(_02140_),
    .S1(_02135_),
    .X(_06011_));
 sky130_fd_sc_hd__or2_2 _12224_ (.A(_02139_),
    .B(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__o311a_2 _12225_ (.A1(_02147_),
    .A2(_06008_),
    .A3(_06010_),
    .B1(_02129_),
    .C1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__or3_2 _12226_ (.A(_00004_),
    .B(_06006_),
    .C(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__buf_1 _12227_ (.A(_02149_),
    .X(_06015_));
 sky130_fd_sc_hd__mux4_2 _12228_ (.A0(\core.cpuregs[16][5] ),
    .A1(\core.cpuregs[17][5] ),
    .A2(\core.cpuregs[18][5] ),
    .A3(\core.cpuregs[19][5] ),
    .S0(_06015_),
    .S1(_02159_),
    .X(_06016_));
 sky130_fd_sc_hd__nor2_2 _12229_ (.A(_02143_),
    .B(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__buf_1 _12230_ (.A(_02149_),
    .X(_06018_));
 sky130_fd_sc_hd__mux2_2 _12231_ (.A0(\core.cpuregs[20][5] ),
    .A1(\core.cpuregs[21][5] ),
    .S(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__buf_1 _12232_ (.A(_02159_),
    .X(_06020_));
 sky130_fd_sc_hd__mux2_2 _12233_ (.A0(\core.cpuregs[22][5] ),
    .A1(\core.cpuregs[23][5] ),
    .S(_02149_),
    .X(_06021_));
 sky130_fd_sc_hd__a21o_2 _12234_ (.A1(_06020_),
    .A2(_06021_),
    .B1(_02147_),
    .X(_06022_));
 sky130_fd_sc_hd__a21oi_2 _12235_ (.A1(_02167_),
    .A2(_06019_),
    .B1(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__buf_1 _12236_ (.A(_02167_),
    .X(_06024_));
 sky130_fd_sc_hd__buf_1 _12237_ (.A(_06000_),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_2 _12238_ (.A0(\core.cpuregs[28][5] ),
    .A1(\core.cpuregs[29][5] ),
    .S(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__buf_1 _12239_ (.A(_02159_),
    .X(_06027_));
 sky130_fd_sc_hd__mux2_2 _12240_ (.A0(\core.cpuregs[30][5] ),
    .A1(\core.cpuregs[31][5] ),
    .S(_06000_),
    .X(_06028_));
 sky130_fd_sc_hd__a21o_2 _12241_ (.A1(_06027_),
    .A2(_06028_),
    .B1(_02147_),
    .X(_06029_));
 sky130_fd_sc_hd__a21oi_2 _12242_ (.A1(_06024_),
    .A2(_06026_),
    .B1(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__buf_1 _12243_ (.A(_02143_),
    .X(_06031_));
 sky130_fd_sc_hd__mux4_2 _12244_ (.A0(\core.cpuregs[24][5] ),
    .A1(\core.cpuregs[25][5] ),
    .A2(\core.cpuregs[26][5] ),
    .A3(\core.cpuregs[27][5] ),
    .S0(_06015_),
    .S1(_06020_),
    .X(_06032_));
 sky130_fd_sc_hd__o21ai_2 _12245_ (.A1(_06031_),
    .A2(_06032_),
    .B1(_02152_),
    .Y(_06033_));
 sky130_fd_sc_hd__o32a_2 _12246_ (.A1(_02152_),
    .A2(_06017_),
    .A3(_06023_),
    .B1(_06030_),
    .B2(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__nand2_2 _12247_ (.A(_02127_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__or2_2 _12248_ (.A(\core.is_lui_auipc_jal ),
    .B(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .X(_06036_));
 sky130_fd_sc_hd__buf_1 _12249_ (.A(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__a32o_2 _12250_ (.A1(_05998_),
    .A2(_06014_),
    .A3(_06035_),
    .B1(_06037_),
    .B2(\core.decoded_imm[5] ),
    .X(_06038_));
 sky130_fd_sc_hd__mux2_2 _12251_ (.A0(\core.mem_la_wdata[5] ),
    .A1(_06038_),
    .S(_05986_),
    .X(_06039_));
 sky130_fd_sc_hd__buf_1 _12252_ (.A(_06039_),
    .X(_00609_));
 sky130_fd_sc_hd__buf_1 _12253_ (.A(_05987_),
    .X(_06040_));
 sky130_fd_sc_hd__buf_1 _12254_ (.A(_02127_),
    .X(_06041_));
 sky130_fd_sc_hd__buf_1 _12255_ (.A(_02147_),
    .X(_06042_));
 sky130_fd_sc_hd__buf_1 _12256_ (.A(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__buf_1 _12257_ (.A(_06000_),
    .X(_06044_));
 sky130_fd_sc_hd__buf_1 _12258_ (.A(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__buf_1 _12259_ (.A(_06027_),
    .X(_06046_));
 sky130_fd_sc_hd__mux4_2 _12260_ (.A0(\core.cpuregs[12][6] ),
    .A1(\core.cpuregs[13][6] ),
    .A2(\core.cpuregs[14][6] ),
    .A3(\core.cpuregs[15][6] ),
    .S0(_06045_),
    .S1(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__buf_1 _12261_ (.A(_06024_),
    .X(_06048_));
 sky130_fd_sc_hd__buf_1 _12262_ (.A(_06025_),
    .X(_06049_));
 sky130_fd_sc_hd__mux2_2 _12263_ (.A0(\core.cpuregs[8][6] ),
    .A1(\core.cpuregs[9][6] ),
    .S(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_1 _12264_ (.A(_06027_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _12265_ (.A(_06000_),
    .X(_06052_));
 sky130_fd_sc_hd__mux2_2 _12266_ (.A0(\core.cpuregs[10][6] ),
    .A1(\core.cpuregs[11][6] ),
    .S(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__buf_1 _12267_ (.A(_02143_),
    .X(_06054_));
 sky130_fd_sc_hd__a21o_2 _12268_ (.A1(_06051_),
    .A2(_06053_),
    .B1(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__a21o_2 _12269_ (.A1(_06048_),
    .A2(_06050_),
    .B1(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__buf_1 _12270_ (.A(_02152_),
    .X(_06057_));
 sky130_fd_sc_hd__buf_1 _12271_ (.A(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__o211a_2 _12272_ (.A1(_06043_),
    .A2(_06047_),
    .B1(_06056_),
    .C1(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__buf_1 _12273_ (.A(_06042_),
    .X(_06060_));
 sky130_fd_sc_hd__buf_1 _12274_ (.A(_02167_),
    .X(_06061_));
 sky130_fd_sc_hd__buf_1 _12275_ (.A(_06018_),
    .X(_06062_));
 sky130_fd_sc_hd__mux2_2 _12276_ (.A0(\core.cpuregs[4][6] ),
    .A1(\core.cpuregs[5][6] ),
    .S(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__and2_2 _12277_ (.A(_06061_),
    .B(_06063_),
    .X(_06064_));
 sky130_fd_sc_hd__buf_1 _12278_ (.A(_06020_),
    .X(_06065_));
 sky130_fd_sc_hd__buf_1 _12279_ (.A(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__buf_1 _12280_ (.A(_06018_),
    .X(_06067_));
 sky130_fd_sc_hd__mux2_2 _12281_ (.A0(\core.cpuregs[6][6] ),
    .A1(\core.cpuregs[7][6] ),
    .S(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__and2_2 _12282_ (.A(_06066_),
    .B(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__buf_1 _12283_ (.A(_02129_),
    .X(_06070_));
 sky130_fd_sc_hd__buf_1 _12284_ (.A(_02143_),
    .X(_06071_));
 sky130_fd_sc_hd__buf_1 _12285_ (.A(_06015_),
    .X(_06072_));
 sky130_fd_sc_hd__buf_1 _12286_ (.A(_06020_),
    .X(_06073_));
 sky130_fd_sc_hd__mux4_2 _12287_ (.A0(\core.cpuregs[0][6] ),
    .A1(\core.cpuregs[1][6] ),
    .A2(\core.cpuregs[2][6] ),
    .A3(\core.cpuregs[3][6] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__or2_2 _12288_ (.A(_06071_),
    .B(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o311a_2 _12289_ (.A1(_06060_),
    .A2(_06064_),
    .A3(_06069_),
    .B1(_06070_),
    .C1(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__buf_1 _12290_ (.A(_02127_),
    .X(_06077_));
 sky130_fd_sc_hd__buf_1 _12291_ (.A(_02152_),
    .X(_06078_));
 sky130_fd_sc_hd__buf_1 _12292_ (.A(_06031_),
    .X(_06079_));
 sky130_fd_sc_hd__buf_1 _12293_ (.A(_06015_),
    .X(_06080_));
 sky130_fd_sc_hd__mux4_2 _12294_ (.A0(\core.cpuregs[16][6] ),
    .A1(\core.cpuregs[17][6] ),
    .A2(\core.cpuregs[18][6] ),
    .A3(\core.cpuregs[19][6] ),
    .S0(_06080_),
    .S1(_06065_),
    .X(_06081_));
 sky130_fd_sc_hd__nor2_2 _12295_ (.A(_06079_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__buf_1 _12296_ (.A(_02167_),
    .X(_06083_));
 sky130_fd_sc_hd__buf_1 _12297_ (.A(_06018_),
    .X(_06084_));
 sky130_fd_sc_hd__mux2_2 _12298_ (.A0(\core.cpuregs[20][6] ),
    .A1(\core.cpuregs[21][6] ),
    .S(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__buf_1 _12299_ (.A(_06027_),
    .X(_06086_));
 sky130_fd_sc_hd__mux2_2 _12300_ (.A0(\core.cpuregs[22][6] ),
    .A1(\core.cpuregs[23][6] ),
    .S(_06025_),
    .X(_06087_));
 sky130_fd_sc_hd__buf_1 _12301_ (.A(_02147_),
    .X(_06088_));
 sky130_fd_sc_hd__a21o_2 _12302_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__a21oi_2 _12303_ (.A1(_06083_),
    .A2(_06085_),
    .B1(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__buf_1 _12304_ (.A(_06024_),
    .X(_06091_));
 sky130_fd_sc_hd__buf_1 _12305_ (.A(_06052_),
    .X(_06092_));
 sky130_fd_sc_hd__mux2_2 _12306_ (.A0(\core.cpuregs[28][6] ),
    .A1(\core.cpuregs[29][6] ),
    .S(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__buf_1 _12307_ (.A(_06027_),
    .X(_06094_));
 sky130_fd_sc_hd__mux2_2 _12308_ (.A0(\core.cpuregs[30][6] ),
    .A1(\core.cpuregs[31][6] ),
    .S(_06044_),
    .X(_06095_));
 sky130_fd_sc_hd__a21o_2 _12309_ (.A1(_06094_),
    .A2(_06095_),
    .B1(_06042_),
    .X(_06096_));
 sky130_fd_sc_hd__a21oi_2 _12310_ (.A1(_06091_),
    .A2(_06093_),
    .B1(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__buf_1 _12311_ (.A(_02143_),
    .X(_06098_));
 sky130_fd_sc_hd__buf_1 _12312_ (.A(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__buf_1 _12313_ (.A(_06018_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_1 _12314_ (.A(_06020_),
    .X(_06101_));
 sky130_fd_sc_hd__mux4_2 _12315_ (.A0(\core.cpuregs[24][6] ),
    .A1(\core.cpuregs[25][6] ),
    .A2(\core.cpuregs[26][6] ),
    .A3(\core.cpuregs[27][6] ),
    .S0(_06100_),
    .S1(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__buf_1 _12316_ (.A(_02152_),
    .X(_06103_));
 sky130_fd_sc_hd__o21ai_2 _12317_ (.A1(_06099_),
    .A2(_06102_),
    .B1(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__o32a_2 _12318_ (.A1(_06078_),
    .A2(_06082_),
    .A3(_06090_),
    .B1(_06097_),
    .B2(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nand2_2 _12319_ (.A(_06077_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__buf_1 _12320_ (.A(_05998_),
    .X(_06107_));
 sky130_fd_sc_hd__o311a_2 _12321_ (.A1(_06041_),
    .A2(_06059_),
    .A3(_06076_),
    .B1(_06106_),
    .C1(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__buf_1 _12322_ (.A(_06037_),
    .X(_06109_));
 sky130_fd_sc_hd__nand2_2 _12323_ (.A(_02024_),
    .B(\core.cpu_state[2] ),
    .Y(_06110_));
 sky130_fd_sc_hd__buf_1 _12324_ (.A(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__a21o_2 _12325_ (.A1(\core.decoded_imm[6] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__o22a_2 _12326_ (.A1(\core.mem_la_wdata[6] ),
    .A2(_06040_),
    .B1(_06108_),
    .B2(_06112_),
    .X(_00610_));
 sky130_fd_sc_hd__mux4_2 _12327_ (.A0(\core.cpuregs[12][7] ),
    .A1(\core.cpuregs[13][7] ),
    .A2(\core.cpuregs[14][7] ),
    .A3(\core.cpuregs[15][7] ),
    .S0(_06045_),
    .S1(_06046_),
    .X(_06113_));
 sky130_fd_sc_hd__mux2_2 _12328_ (.A0(\core.cpuregs[8][7] ),
    .A1(\core.cpuregs[9][7] ),
    .S(_06049_),
    .X(_06114_));
 sky130_fd_sc_hd__mux2_2 _12329_ (.A0(\core.cpuregs[10][7] ),
    .A1(\core.cpuregs[11][7] ),
    .S(_06052_),
    .X(_06115_));
 sky130_fd_sc_hd__a21o_2 _12330_ (.A1(_06051_),
    .A2(_06115_),
    .B1(_06054_),
    .X(_06116_));
 sky130_fd_sc_hd__a21o_2 _12331_ (.A1(_06048_),
    .A2(_06114_),
    .B1(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__o211a_2 _12332_ (.A1(_06043_),
    .A2(_06113_),
    .B1(_06117_),
    .C1(_06058_),
    .X(_06118_));
 sky130_fd_sc_hd__mux2_2 _12333_ (.A0(\core.cpuregs[4][7] ),
    .A1(\core.cpuregs[5][7] ),
    .S(_06062_),
    .X(_06119_));
 sky130_fd_sc_hd__and2_2 _12334_ (.A(_06061_),
    .B(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__mux2_2 _12335_ (.A0(\core.cpuregs[6][7] ),
    .A1(\core.cpuregs[7][7] ),
    .S(_06067_),
    .X(_06121_));
 sky130_fd_sc_hd__and2_2 _12336_ (.A(_06066_),
    .B(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__mux4_2 _12337_ (.A0(\core.cpuregs[0][7] ),
    .A1(\core.cpuregs[1][7] ),
    .A2(\core.cpuregs[2][7] ),
    .A3(\core.cpuregs[3][7] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06123_));
 sky130_fd_sc_hd__or2_2 _12338_ (.A(_06071_),
    .B(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__o311a_2 _12339_ (.A1(_06060_),
    .A2(_06120_),
    .A3(_06122_),
    .B1(_06070_),
    .C1(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__mux4_2 _12340_ (.A0(\core.cpuregs[16][7] ),
    .A1(\core.cpuregs[17][7] ),
    .A2(\core.cpuregs[18][7] ),
    .A3(\core.cpuregs[19][7] ),
    .S0(_06080_),
    .S1(_06065_),
    .X(_06126_));
 sky130_fd_sc_hd__nor2_2 _12341_ (.A(_06079_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__mux2_2 _12342_ (.A0(\core.cpuregs[20][7] ),
    .A1(\core.cpuregs[21][7] ),
    .S(_06084_),
    .X(_06128_));
 sky130_fd_sc_hd__mux2_2 _12343_ (.A0(\core.cpuregs[22][7] ),
    .A1(\core.cpuregs[23][7] ),
    .S(_06025_),
    .X(_06129_));
 sky130_fd_sc_hd__a21o_2 _12344_ (.A1(_06086_),
    .A2(_06129_),
    .B1(_06088_),
    .X(_06130_));
 sky130_fd_sc_hd__a21oi_2 _12345_ (.A1(_06083_),
    .A2(_06128_),
    .B1(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__mux2_2 _12346_ (.A0(\core.cpuregs[28][7] ),
    .A1(\core.cpuregs[29][7] ),
    .S(_06092_),
    .X(_06132_));
 sky130_fd_sc_hd__mux2_2 _12347_ (.A0(\core.cpuregs[30][7] ),
    .A1(\core.cpuregs[31][7] ),
    .S(_06044_),
    .X(_06133_));
 sky130_fd_sc_hd__a21o_2 _12348_ (.A1(_06094_),
    .A2(_06133_),
    .B1(_06042_),
    .X(_06134_));
 sky130_fd_sc_hd__a21oi_2 _12349_ (.A1(_06091_),
    .A2(_06132_),
    .B1(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__mux4_2 _12350_ (.A0(\core.cpuregs[24][7] ),
    .A1(\core.cpuregs[25][7] ),
    .A2(\core.cpuregs[26][7] ),
    .A3(\core.cpuregs[27][7] ),
    .S0(_06100_),
    .S1(_06101_),
    .X(_06136_));
 sky130_fd_sc_hd__o21ai_2 _12351_ (.A1(_06099_),
    .A2(_06136_),
    .B1(_06103_),
    .Y(_06137_));
 sky130_fd_sc_hd__o32a_2 _12352_ (.A1(_06078_),
    .A2(_06127_),
    .A3(_06131_),
    .B1(_06135_),
    .B2(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__nand2_2 _12353_ (.A(_06077_),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__o311a_2 _12354_ (.A1(_06041_),
    .A2(_06118_),
    .A3(_06125_),
    .B1(_06139_),
    .C1(_06107_),
    .X(_06140_));
 sky130_fd_sc_hd__a21o_2 _12355_ (.A1(\core.decoded_imm[7] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06141_));
 sky130_fd_sc_hd__o22a_2 _12356_ (.A1(\core.mem_la_wdata[7] ),
    .A2(_06040_),
    .B1(_06140_),
    .B2(_06141_),
    .X(_00611_));
 sky130_fd_sc_hd__mux4_2 _12357_ (.A0(\core.cpuregs[12][8] ),
    .A1(\core.cpuregs[13][8] ),
    .A2(\core.cpuregs[14][8] ),
    .A3(\core.cpuregs[15][8] ),
    .S0(_06045_),
    .S1(_06046_),
    .X(_06142_));
 sky130_fd_sc_hd__mux2_2 _12358_ (.A0(\core.cpuregs[8][8] ),
    .A1(\core.cpuregs[9][8] ),
    .S(_06049_),
    .X(_06143_));
 sky130_fd_sc_hd__buf_1 _12359_ (.A(_06027_),
    .X(_06144_));
 sky130_fd_sc_hd__mux2_2 _12360_ (.A0(\core.cpuregs[10][8] ),
    .A1(\core.cpuregs[11][8] ),
    .S(_06052_),
    .X(_06145_));
 sky130_fd_sc_hd__a21o_2 _12361_ (.A1(_06144_),
    .A2(_06145_),
    .B1(_06054_),
    .X(_06146_));
 sky130_fd_sc_hd__a21o_2 _12362_ (.A1(_06048_),
    .A2(_06143_),
    .B1(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__o211a_2 _12363_ (.A1(_06043_),
    .A2(_06142_),
    .B1(_06147_),
    .C1(_06058_),
    .X(_06148_));
 sky130_fd_sc_hd__buf_1 _12364_ (.A(_02167_),
    .X(_06149_));
 sky130_fd_sc_hd__mux2_2 _12365_ (.A0(\core.cpuregs[4][8] ),
    .A1(\core.cpuregs[5][8] ),
    .S(_06062_),
    .X(_06150_));
 sky130_fd_sc_hd__and2_2 _12366_ (.A(_06149_),
    .B(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__mux2_2 _12367_ (.A0(\core.cpuregs[6][8] ),
    .A1(\core.cpuregs[7][8] ),
    .S(_06067_),
    .X(_06152_));
 sky130_fd_sc_hd__and2_2 _12368_ (.A(_06066_),
    .B(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__buf_1 _12369_ (.A(_06015_),
    .X(_06154_));
 sky130_fd_sc_hd__mux4_2 _12370_ (.A0(\core.cpuregs[0][8] ),
    .A1(\core.cpuregs[1][8] ),
    .A2(\core.cpuregs[2][8] ),
    .A3(\core.cpuregs[3][8] ),
    .S0(_06154_),
    .S1(_06073_),
    .X(_06155_));
 sky130_fd_sc_hd__or2_2 _12371_ (.A(_06071_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__o311a_2 _12372_ (.A1(_06060_),
    .A2(_06151_),
    .A3(_06153_),
    .B1(_06070_),
    .C1(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__buf_1 _12373_ (.A(_06020_),
    .X(_06158_));
 sky130_fd_sc_hd__mux4_2 _12374_ (.A0(\core.cpuregs[16][8] ),
    .A1(\core.cpuregs[17][8] ),
    .A2(\core.cpuregs[18][8] ),
    .A3(\core.cpuregs[19][8] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__nor2_2 _12375_ (.A(_06079_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__buf_1 _12376_ (.A(_06018_),
    .X(_06161_));
 sky130_fd_sc_hd__mux2_2 _12377_ (.A0(\core.cpuregs[20][8] ),
    .A1(\core.cpuregs[21][8] ),
    .S(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__mux2_2 _12378_ (.A0(\core.cpuregs[22][8] ),
    .A1(\core.cpuregs[23][8] ),
    .S(_06025_),
    .X(_06163_));
 sky130_fd_sc_hd__a21o_2 _12379_ (.A1(_06086_),
    .A2(_06163_),
    .B1(_06088_),
    .X(_06164_));
 sky130_fd_sc_hd__a21oi_2 _12380_ (.A1(_06083_),
    .A2(_06162_),
    .B1(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__mux2_2 _12381_ (.A0(\core.cpuregs[28][8] ),
    .A1(\core.cpuregs[29][8] ),
    .S(_06092_),
    .X(_06166_));
 sky130_fd_sc_hd__mux2_2 _12382_ (.A0(\core.cpuregs[30][8] ),
    .A1(\core.cpuregs[31][8] ),
    .S(_06044_),
    .X(_06167_));
 sky130_fd_sc_hd__a21o_2 _12383_ (.A1(_06094_),
    .A2(_06167_),
    .B1(_06042_),
    .X(_06168_));
 sky130_fd_sc_hd__a21oi_2 _12384_ (.A1(_06091_),
    .A2(_06166_),
    .B1(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__mux4_2 _12385_ (.A0(\core.cpuregs[24][8] ),
    .A1(\core.cpuregs[25][8] ),
    .A2(\core.cpuregs[26][8] ),
    .A3(\core.cpuregs[27][8] ),
    .S0(_06100_),
    .S1(_06101_),
    .X(_06170_));
 sky130_fd_sc_hd__o21ai_2 _12386_ (.A1(_06099_),
    .A2(_06170_),
    .B1(_06103_),
    .Y(_06171_));
 sky130_fd_sc_hd__o32a_2 _12387_ (.A1(_06078_),
    .A2(_06160_),
    .A3(_06165_),
    .B1(_06169_),
    .B2(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__nand2_2 _12388_ (.A(_06077_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__o311a_2 _12389_ (.A1(_06041_),
    .A2(_06148_),
    .A3(_06157_),
    .B1(_06173_),
    .C1(_06107_),
    .X(_06174_));
 sky130_fd_sc_hd__a21o_2 _12390_ (.A1(\core.decoded_imm[8] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06175_));
 sky130_fd_sc_hd__o22a_2 _12391_ (.A1(\core.pcpi_rs2[8] ),
    .A2(_06040_),
    .B1(_06174_),
    .B2(_06175_),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_2 _12392_ (.A0(\core.cpuregs[12][9] ),
    .A1(\core.cpuregs[13][9] ),
    .A2(\core.cpuregs[14][9] ),
    .A3(\core.cpuregs[15][9] ),
    .S0(_06045_),
    .S1(_06046_),
    .X(_06176_));
 sky130_fd_sc_hd__mux2_2 _12393_ (.A0(\core.cpuregs[8][9] ),
    .A1(\core.cpuregs[9][9] ),
    .S(_06049_),
    .X(_06177_));
 sky130_fd_sc_hd__mux2_2 _12394_ (.A0(\core.cpuregs[10][9] ),
    .A1(\core.cpuregs[11][9] ),
    .S(_06052_),
    .X(_06178_));
 sky130_fd_sc_hd__a21o_2 _12395_ (.A1(_06144_),
    .A2(_06178_),
    .B1(_06054_),
    .X(_06179_));
 sky130_fd_sc_hd__a21o_2 _12396_ (.A1(_06048_),
    .A2(_06177_),
    .B1(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__o211a_2 _12397_ (.A1(_06043_),
    .A2(_06176_),
    .B1(_06180_),
    .C1(_06058_),
    .X(_06181_));
 sky130_fd_sc_hd__mux2_2 _12398_ (.A0(\core.cpuregs[4][9] ),
    .A1(\core.cpuregs[5][9] ),
    .S(_06062_),
    .X(_06182_));
 sky130_fd_sc_hd__and2_2 _12399_ (.A(_06149_),
    .B(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__mux2_2 _12400_ (.A0(\core.cpuregs[6][9] ),
    .A1(\core.cpuregs[7][9] ),
    .S(_06067_),
    .X(_06184_));
 sky130_fd_sc_hd__and2_2 _12401_ (.A(_06066_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__mux4_2 _12402_ (.A0(\core.cpuregs[0][9] ),
    .A1(\core.cpuregs[1][9] ),
    .A2(\core.cpuregs[2][9] ),
    .A3(\core.cpuregs[3][9] ),
    .S0(_06154_),
    .S1(_06073_),
    .X(_06186_));
 sky130_fd_sc_hd__or2_2 _12403_ (.A(_06071_),
    .B(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__o311a_2 _12404_ (.A1(_06060_),
    .A2(_06183_),
    .A3(_06185_),
    .B1(_06070_),
    .C1(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__mux4_2 _12405_ (.A0(\core.cpuregs[16][9] ),
    .A1(\core.cpuregs[17][9] ),
    .A2(\core.cpuregs[18][9] ),
    .A3(\core.cpuregs[19][9] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06189_));
 sky130_fd_sc_hd__nor2_2 _12406_ (.A(_06079_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__mux2_2 _12407_ (.A0(\core.cpuregs[20][9] ),
    .A1(\core.cpuregs[21][9] ),
    .S(_06161_),
    .X(_06191_));
 sky130_fd_sc_hd__mux2_2 _12408_ (.A0(\core.cpuregs[22][9] ),
    .A1(\core.cpuregs[23][9] ),
    .S(_06025_),
    .X(_06192_));
 sky130_fd_sc_hd__a21o_2 _12409_ (.A1(_06086_),
    .A2(_06192_),
    .B1(_06088_),
    .X(_06193_));
 sky130_fd_sc_hd__a21oi_2 _12410_ (.A1(_06083_),
    .A2(_06191_),
    .B1(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__mux2_2 _12411_ (.A0(\core.cpuregs[28][9] ),
    .A1(\core.cpuregs[29][9] ),
    .S(_06092_),
    .X(_06195_));
 sky130_fd_sc_hd__mux2_2 _12412_ (.A0(\core.cpuregs[30][9] ),
    .A1(\core.cpuregs[31][9] ),
    .S(_06044_),
    .X(_06196_));
 sky130_fd_sc_hd__buf_1 _12413_ (.A(_02147_),
    .X(_06197_));
 sky130_fd_sc_hd__a21o_2 _12414_ (.A1(_06094_),
    .A2(_06196_),
    .B1(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__a21oi_2 _12415_ (.A1(_06091_),
    .A2(_06195_),
    .B1(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__mux4_2 _12416_ (.A0(\core.cpuregs[24][9] ),
    .A1(\core.cpuregs[25][9] ),
    .A2(\core.cpuregs[26][9] ),
    .A3(\core.cpuregs[27][9] ),
    .S0(_06100_),
    .S1(_06101_),
    .X(_06200_));
 sky130_fd_sc_hd__o21ai_2 _12417_ (.A1(_06099_),
    .A2(_06200_),
    .B1(_06103_),
    .Y(_06201_));
 sky130_fd_sc_hd__o32a_2 _12418_ (.A1(_06078_),
    .A2(_06190_),
    .A3(_06194_),
    .B1(_06199_),
    .B2(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__nand2_2 _12419_ (.A(_06077_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__o311a_2 _12420_ (.A1(_06041_),
    .A2(_06181_),
    .A3(_06188_),
    .B1(_06203_),
    .C1(_06107_),
    .X(_06204_));
 sky130_fd_sc_hd__a21o_2 _12421_ (.A1(\core.decoded_imm[9] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06205_));
 sky130_fd_sc_hd__o22a_2 _12422_ (.A1(\core.pcpi_rs2[9] ),
    .A2(_06040_),
    .B1(_06204_),
    .B2(_06205_),
    .X(_00613_));
 sky130_fd_sc_hd__buf_1 _12423_ (.A(_06027_),
    .X(_06206_));
 sky130_fd_sc_hd__mux4_2 _12424_ (.A0(\core.cpuregs[12][10] ),
    .A1(\core.cpuregs[13][10] ),
    .A2(\core.cpuregs[14][10] ),
    .A3(\core.cpuregs[15][10] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__buf_1 _12425_ (.A(_06024_),
    .X(_06208_));
 sky130_fd_sc_hd__mux2_2 _12426_ (.A0(\core.cpuregs[8][10] ),
    .A1(\core.cpuregs[9][10] ),
    .S(_06049_),
    .X(_06209_));
 sky130_fd_sc_hd__mux2_2 _12427_ (.A0(\core.cpuregs[10][10] ),
    .A1(\core.cpuregs[11][10] ),
    .S(_06052_),
    .X(_06210_));
 sky130_fd_sc_hd__a21o_2 _12428_ (.A1(_06144_),
    .A2(_06210_),
    .B1(_06054_),
    .X(_06211_));
 sky130_fd_sc_hd__a21o_2 _12429_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__o211a_2 _12430_ (.A1(_06043_),
    .A2(_06207_),
    .B1(_06212_),
    .C1(_06058_),
    .X(_06213_));
 sky130_fd_sc_hd__buf_1 _12431_ (.A(_06042_),
    .X(_06214_));
 sky130_fd_sc_hd__mux2_2 _12432_ (.A0(\core.cpuregs[4][10] ),
    .A1(\core.cpuregs[5][10] ),
    .S(_06062_),
    .X(_06215_));
 sky130_fd_sc_hd__and2_2 _12433_ (.A(_06149_),
    .B(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__mux2_2 _12434_ (.A0(\core.cpuregs[6][10] ),
    .A1(\core.cpuregs[7][10] ),
    .S(_06067_),
    .X(_06217_));
 sky130_fd_sc_hd__and2_2 _12435_ (.A(_06066_),
    .B(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__mux4_2 _12436_ (.A0(\core.cpuregs[0][10] ),
    .A1(\core.cpuregs[1][10] ),
    .A2(\core.cpuregs[2][10] ),
    .A3(\core.cpuregs[3][10] ),
    .S0(_06154_),
    .S1(_06073_),
    .X(_06219_));
 sky130_fd_sc_hd__or2_2 _12437_ (.A(_06071_),
    .B(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__o311a_2 _12438_ (.A1(_06214_),
    .A2(_06216_),
    .A3(_06218_),
    .B1(_06070_),
    .C1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__buf_1 _12439_ (.A(_02127_),
    .X(_06222_));
 sky130_fd_sc_hd__buf_1 _12440_ (.A(_02152_),
    .X(_06223_));
 sky130_fd_sc_hd__buf_1 _12441_ (.A(_06031_),
    .X(_06224_));
 sky130_fd_sc_hd__mux4_2 _12442_ (.A0(\core.cpuregs[16][10] ),
    .A1(\core.cpuregs[17][10] ),
    .A2(\core.cpuregs[18][10] ),
    .A3(\core.cpuregs[19][10] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_2 _12443_ (.A(_06224_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__mux2_2 _12444_ (.A0(\core.cpuregs[20][10] ),
    .A1(\core.cpuregs[21][10] ),
    .S(_06161_),
    .X(_06227_));
 sky130_fd_sc_hd__mux2_2 _12445_ (.A0(\core.cpuregs[22][10] ),
    .A1(\core.cpuregs[23][10] ),
    .S(_06025_),
    .X(_06228_));
 sky130_fd_sc_hd__a21o_2 _12446_ (.A1(_06086_),
    .A2(_06228_),
    .B1(_06088_),
    .X(_06229_));
 sky130_fd_sc_hd__a21oi_2 _12447_ (.A1(_06083_),
    .A2(_06227_),
    .B1(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__buf_1 _12448_ (.A(_06052_),
    .X(_06231_));
 sky130_fd_sc_hd__mux2_2 _12449_ (.A0(\core.cpuregs[28][10] ),
    .A1(\core.cpuregs[29][10] ),
    .S(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__buf_1 _12450_ (.A(_06015_),
    .X(_06233_));
 sky130_fd_sc_hd__mux2_2 _12451_ (.A0(\core.cpuregs[30][10] ),
    .A1(\core.cpuregs[31][10] ),
    .S(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__a21o_2 _12452_ (.A1(_06094_),
    .A2(_06234_),
    .B1(_06197_),
    .X(_06235_));
 sky130_fd_sc_hd__a21oi_2 _12453_ (.A1(_06091_),
    .A2(_06232_),
    .B1(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__buf_1 _12454_ (.A(_06015_),
    .X(_06237_));
 sky130_fd_sc_hd__mux4_2 _12455_ (.A0(\core.cpuregs[24][10] ),
    .A1(\core.cpuregs[25][10] ),
    .A2(\core.cpuregs[26][10] ),
    .A3(\core.cpuregs[27][10] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06238_));
 sky130_fd_sc_hd__o21ai_2 _12456_ (.A1(_06099_),
    .A2(_06238_),
    .B1(_06103_),
    .Y(_06239_));
 sky130_fd_sc_hd__o32a_2 _12457_ (.A1(_06223_),
    .A2(_06226_),
    .A3(_06230_),
    .B1(_06236_),
    .B2(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__nand2_2 _12458_ (.A(_06222_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__o311a_2 _12459_ (.A1(_06041_),
    .A2(_06213_),
    .A3(_06221_),
    .B1(_06241_),
    .C1(_06107_),
    .X(_06242_));
 sky130_fd_sc_hd__a21o_2 _12460_ (.A1(\core.decoded_imm[10] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06243_));
 sky130_fd_sc_hd__o22a_2 _12461_ (.A1(\core.pcpi_rs2[10] ),
    .A2(_06040_),
    .B1(_06242_),
    .B2(_06243_),
    .X(_00614_));
 sky130_fd_sc_hd__mux4_2 _12462_ (.A0(\core.cpuregs[12][11] ),
    .A1(\core.cpuregs[13][11] ),
    .A2(\core.cpuregs[14][11] ),
    .A3(\core.cpuregs[15][11] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06244_));
 sky130_fd_sc_hd__mux2_2 _12463_ (.A0(\core.cpuregs[8][11] ),
    .A1(\core.cpuregs[9][11] ),
    .S(_06049_),
    .X(_06245_));
 sky130_fd_sc_hd__buf_1 _12464_ (.A(_06000_),
    .X(_06246_));
 sky130_fd_sc_hd__mux2_2 _12465_ (.A0(\core.cpuregs[10][11] ),
    .A1(\core.cpuregs[11][11] ),
    .S(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a21o_2 _12466_ (.A1(_06144_),
    .A2(_06247_),
    .B1(_06054_),
    .X(_06248_));
 sky130_fd_sc_hd__a21o_2 _12467_ (.A1(_06208_),
    .A2(_06245_),
    .B1(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__o211a_2 _12468_ (.A1(_06043_),
    .A2(_06244_),
    .B1(_06249_),
    .C1(_06058_),
    .X(_06250_));
 sky130_fd_sc_hd__mux2_2 _12469_ (.A0(\core.cpuregs[4][11] ),
    .A1(\core.cpuregs[5][11] ),
    .S(_06062_),
    .X(_06251_));
 sky130_fd_sc_hd__and2_2 _12470_ (.A(_06149_),
    .B(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__mux2_2 _12471_ (.A0(\core.cpuregs[6][11] ),
    .A1(\core.cpuregs[7][11] ),
    .S(_06067_),
    .X(_06253_));
 sky130_fd_sc_hd__and2_2 _12472_ (.A(_06066_),
    .B(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__mux4_2 _12473_ (.A0(\core.cpuregs[0][11] ),
    .A1(\core.cpuregs[1][11] ),
    .A2(\core.cpuregs[2][11] ),
    .A3(\core.cpuregs[3][11] ),
    .S0(_06154_),
    .S1(_06073_),
    .X(_06255_));
 sky130_fd_sc_hd__or2_2 _12474_ (.A(_06071_),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__o311a_2 _12475_ (.A1(_06214_),
    .A2(_06252_),
    .A3(_06254_),
    .B1(_06070_),
    .C1(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__mux4_2 _12476_ (.A0(\core.cpuregs[16][11] ),
    .A1(\core.cpuregs[17][11] ),
    .A2(\core.cpuregs[18][11] ),
    .A3(\core.cpuregs[19][11] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06258_));
 sky130_fd_sc_hd__nor2_2 _12477_ (.A(_06224_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__mux2_2 _12478_ (.A0(\core.cpuregs[20][11] ),
    .A1(\core.cpuregs[21][11] ),
    .S(_06161_),
    .X(_06260_));
 sky130_fd_sc_hd__mux2_2 _12479_ (.A0(\core.cpuregs[22][11] ),
    .A1(\core.cpuregs[23][11] ),
    .S(_06025_),
    .X(_06261_));
 sky130_fd_sc_hd__a21o_2 _12480_ (.A1(_06086_),
    .A2(_06261_),
    .B1(_06088_),
    .X(_06262_));
 sky130_fd_sc_hd__a21oi_2 _12481_ (.A1(_06083_),
    .A2(_06260_),
    .B1(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__mux2_2 _12482_ (.A0(\core.cpuregs[28][11] ),
    .A1(\core.cpuregs[29][11] ),
    .S(_06231_),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_2 _12483_ (.A0(\core.cpuregs[30][11] ),
    .A1(\core.cpuregs[31][11] ),
    .S(_06233_),
    .X(_06265_));
 sky130_fd_sc_hd__a21o_2 _12484_ (.A1(_06094_),
    .A2(_06265_),
    .B1(_06197_),
    .X(_06266_));
 sky130_fd_sc_hd__a21oi_2 _12485_ (.A1(_06091_),
    .A2(_06264_),
    .B1(_06266_),
    .Y(_06267_));
 sky130_fd_sc_hd__mux4_2 _12486_ (.A0(\core.cpuregs[24][11] ),
    .A1(\core.cpuregs[25][11] ),
    .A2(\core.cpuregs[26][11] ),
    .A3(\core.cpuregs[27][11] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06268_));
 sky130_fd_sc_hd__o21ai_2 _12487_ (.A1(_06099_),
    .A2(_06268_),
    .B1(_06103_),
    .Y(_06269_));
 sky130_fd_sc_hd__o32a_2 _12488_ (.A1(_06223_),
    .A2(_06259_),
    .A3(_06263_),
    .B1(_06267_),
    .B2(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__nand2_2 _12489_ (.A(_06222_),
    .B(_06270_),
    .Y(_06271_));
 sky130_fd_sc_hd__o311a_2 _12490_ (.A1(_06041_),
    .A2(_06250_),
    .A3(_06257_),
    .B1(_06271_),
    .C1(_06107_),
    .X(_06272_));
 sky130_fd_sc_hd__a21o_2 _12491_ (.A1(\core.decoded_imm[11] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06273_));
 sky130_fd_sc_hd__o22a_2 _12492_ (.A1(\core.pcpi_rs2[11] ),
    .A2(_06040_),
    .B1(_06272_),
    .B2(_06273_),
    .X(_00615_));
 sky130_fd_sc_hd__mux4_2 _12493_ (.A0(\core.cpuregs[12][12] ),
    .A1(\core.cpuregs[13][12] ),
    .A2(\core.cpuregs[14][12] ),
    .A3(\core.cpuregs[15][12] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06274_));
 sky130_fd_sc_hd__mux2_2 _12494_ (.A0(\core.cpuregs[8][12] ),
    .A1(\core.cpuregs[9][12] ),
    .S(_06049_),
    .X(_06275_));
 sky130_fd_sc_hd__mux2_2 _12495_ (.A0(\core.cpuregs[10][12] ),
    .A1(\core.cpuregs[11][12] ),
    .S(_06246_),
    .X(_06276_));
 sky130_fd_sc_hd__a21o_2 _12496_ (.A1(_06144_),
    .A2(_06276_),
    .B1(_06054_),
    .X(_06277_));
 sky130_fd_sc_hd__a21o_2 _12497_ (.A1(_06208_),
    .A2(_06275_),
    .B1(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__o211a_2 _12498_ (.A1(_06043_),
    .A2(_06274_),
    .B1(_06278_),
    .C1(_06058_),
    .X(_06279_));
 sky130_fd_sc_hd__mux2_2 _12499_ (.A0(\core.cpuregs[4][12] ),
    .A1(\core.cpuregs[5][12] ),
    .S(_06062_),
    .X(_06280_));
 sky130_fd_sc_hd__and2_2 _12500_ (.A(_06149_),
    .B(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__buf_1 _12501_ (.A(_06018_),
    .X(_06282_));
 sky130_fd_sc_hd__mux2_2 _12502_ (.A0(\core.cpuregs[6][12] ),
    .A1(\core.cpuregs[7][12] ),
    .S(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__and2_2 _12503_ (.A(_06066_),
    .B(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__buf_1 _12504_ (.A(_02159_),
    .X(_06285_));
 sky130_fd_sc_hd__mux4_2 _12505_ (.A0(\core.cpuregs[0][12] ),
    .A1(\core.cpuregs[1][12] ),
    .A2(\core.cpuregs[2][12] ),
    .A3(\core.cpuregs[3][12] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06286_));
 sky130_fd_sc_hd__or2_2 _12506_ (.A(_06071_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__o311a_2 _12507_ (.A1(_06214_),
    .A2(_06281_),
    .A3(_06284_),
    .B1(_06070_),
    .C1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__mux4_2 _12508_ (.A0(\core.cpuregs[16][12] ),
    .A1(\core.cpuregs[17][12] ),
    .A2(\core.cpuregs[18][12] ),
    .A3(\core.cpuregs[19][12] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_2 _12509_ (.A(_06224_),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__mux2_2 _12510_ (.A0(\core.cpuregs[20][12] ),
    .A1(\core.cpuregs[21][12] ),
    .S(_06161_),
    .X(_06291_));
 sky130_fd_sc_hd__buf_1 _12511_ (.A(_06020_),
    .X(_06292_));
 sky130_fd_sc_hd__buf_1 _12512_ (.A(_06000_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2_2 _12513_ (.A0(\core.cpuregs[22][12] ),
    .A1(\core.cpuregs[23][12] ),
    .S(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__a21o_2 _12514_ (.A1(_06292_),
    .A2(_06294_),
    .B1(_06088_),
    .X(_06295_));
 sky130_fd_sc_hd__a21oi_2 _12515_ (.A1(_06083_),
    .A2(_06291_),
    .B1(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__mux2_2 _12516_ (.A0(\core.cpuregs[28][12] ),
    .A1(\core.cpuregs[29][12] ),
    .S(_06231_),
    .X(_06297_));
 sky130_fd_sc_hd__mux2_2 _12517_ (.A0(\core.cpuregs[30][12] ),
    .A1(\core.cpuregs[31][12] ),
    .S(_06233_),
    .X(_06298_));
 sky130_fd_sc_hd__a21o_2 _12518_ (.A1(_06094_),
    .A2(_06298_),
    .B1(_06197_),
    .X(_06299_));
 sky130_fd_sc_hd__a21oi_2 _12519_ (.A1(_06091_),
    .A2(_06297_),
    .B1(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__mux4_2 _12520_ (.A0(\core.cpuregs[24][12] ),
    .A1(\core.cpuregs[25][12] ),
    .A2(\core.cpuregs[26][12] ),
    .A3(\core.cpuregs[27][12] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06301_));
 sky130_fd_sc_hd__o21ai_2 _12521_ (.A1(_06099_),
    .A2(_06301_),
    .B1(_06103_),
    .Y(_06302_));
 sky130_fd_sc_hd__o32a_2 _12522_ (.A1(_06223_),
    .A2(_06290_),
    .A3(_06296_),
    .B1(_06300_),
    .B2(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__nand2_2 _12523_ (.A(_06222_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__o311a_2 _12524_ (.A1(_06041_),
    .A2(_06279_),
    .A3(_06288_),
    .B1(_06304_),
    .C1(_06107_),
    .X(_06305_));
 sky130_fd_sc_hd__a21o_2 _12525_ (.A1(\core.decoded_imm[12] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06306_));
 sky130_fd_sc_hd__o22a_2 _12526_ (.A1(\core.pcpi_rs2[12] ),
    .A2(_06040_),
    .B1(_06305_),
    .B2(_06306_),
    .X(_00616_));
 sky130_fd_sc_hd__mux4_2 _12527_ (.A0(\core.cpuregs[12][13] ),
    .A1(\core.cpuregs[13][13] ),
    .A2(\core.cpuregs[14][13] ),
    .A3(\core.cpuregs[15][13] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06307_));
 sky130_fd_sc_hd__mux2_2 _12528_ (.A0(\core.cpuregs[8][13] ),
    .A1(\core.cpuregs[9][13] ),
    .S(_06049_),
    .X(_06308_));
 sky130_fd_sc_hd__mux2_2 _12529_ (.A0(\core.cpuregs[10][13] ),
    .A1(\core.cpuregs[11][13] ),
    .S(_06246_),
    .X(_06309_));
 sky130_fd_sc_hd__a21o_2 _12530_ (.A1(_06144_),
    .A2(_06309_),
    .B1(_06054_),
    .X(_06310_));
 sky130_fd_sc_hd__a21o_2 _12531_ (.A1(_06208_),
    .A2(_06308_),
    .B1(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__o211a_2 _12532_ (.A1(_06043_),
    .A2(_06307_),
    .B1(_06311_),
    .C1(_06058_),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_2 _12533_ (.A0(\core.cpuregs[4][13] ),
    .A1(\core.cpuregs[5][13] ),
    .S(_06062_),
    .X(_06313_));
 sky130_fd_sc_hd__and2_2 _12534_ (.A(_06149_),
    .B(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_2 _12535_ (.A0(\core.cpuregs[6][13] ),
    .A1(\core.cpuregs[7][13] ),
    .S(_06282_),
    .X(_06315_));
 sky130_fd_sc_hd__and2_2 _12536_ (.A(_06066_),
    .B(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__mux4_2 _12537_ (.A0(\core.cpuregs[0][13] ),
    .A1(\core.cpuregs[1][13] ),
    .A2(\core.cpuregs[2][13] ),
    .A3(\core.cpuregs[3][13] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06317_));
 sky130_fd_sc_hd__or2_2 _12538_ (.A(_06071_),
    .B(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__o311a_2 _12539_ (.A1(_06214_),
    .A2(_06314_),
    .A3(_06316_),
    .B1(_06070_),
    .C1(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__mux4_2 _12540_ (.A0(\core.cpuregs[16][13] ),
    .A1(\core.cpuregs[17][13] ),
    .A2(\core.cpuregs[18][13] ),
    .A3(\core.cpuregs[19][13] ),
    .S0(_06080_),
    .S1(_06158_),
    .X(_06320_));
 sky130_fd_sc_hd__nor2_2 _12541_ (.A(_06224_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__mux2_2 _12542_ (.A0(\core.cpuregs[20][13] ),
    .A1(\core.cpuregs[21][13] ),
    .S(_06161_),
    .X(_06322_));
 sky130_fd_sc_hd__mux2_2 _12543_ (.A0(\core.cpuregs[22][13] ),
    .A1(\core.cpuregs[23][13] ),
    .S(_06293_),
    .X(_06323_));
 sky130_fd_sc_hd__buf_1 _12544_ (.A(_02147_),
    .X(_06324_));
 sky130_fd_sc_hd__a21o_2 _12545_ (.A1(_06292_),
    .A2(_06323_),
    .B1(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__a21oi_2 _12546_ (.A1(_06083_),
    .A2(_06322_),
    .B1(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__mux2_2 _12547_ (.A0(\core.cpuregs[28][13] ),
    .A1(\core.cpuregs[29][13] ),
    .S(_06231_),
    .X(_06327_));
 sky130_fd_sc_hd__mux2_2 _12548_ (.A0(\core.cpuregs[30][13] ),
    .A1(\core.cpuregs[31][13] ),
    .S(_06233_),
    .X(_06328_));
 sky130_fd_sc_hd__a21o_2 _12549_ (.A1(_06094_),
    .A2(_06328_),
    .B1(_06197_),
    .X(_06329_));
 sky130_fd_sc_hd__a21oi_2 _12550_ (.A1(_06091_),
    .A2(_06327_),
    .B1(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__mux4_2 _12551_ (.A0(\core.cpuregs[24][13] ),
    .A1(\core.cpuregs[25][13] ),
    .A2(\core.cpuregs[26][13] ),
    .A3(\core.cpuregs[27][13] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06331_));
 sky130_fd_sc_hd__o21ai_2 _12552_ (.A1(_06099_),
    .A2(_06331_),
    .B1(_06103_),
    .Y(_06332_));
 sky130_fd_sc_hd__o32a_2 _12553_ (.A1(_06223_),
    .A2(_06321_),
    .A3(_06326_),
    .B1(_06330_),
    .B2(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__nand2_2 _12554_ (.A(_06222_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__o311a_2 _12555_ (.A1(_06041_),
    .A2(_06312_),
    .A3(_06319_),
    .B1(_06334_),
    .C1(_06107_),
    .X(_06335_));
 sky130_fd_sc_hd__a21o_2 _12556_ (.A1(\core.decoded_imm[13] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06336_));
 sky130_fd_sc_hd__o22a_2 _12557_ (.A1(\core.pcpi_rs2[13] ),
    .A2(_06040_),
    .B1(_06335_),
    .B2(_06336_),
    .X(_00617_));
 sky130_fd_sc_hd__mux4_2 _12558_ (.A0(\core.cpuregs[12][14] ),
    .A1(\core.cpuregs[13][14] ),
    .A2(\core.cpuregs[14][14] ),
    .A3(\core.cpuregs[15][14] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06337_));
 sky130_fd_sc_hd__buf_1 _12559_ (.A(_06025_),
    .X(_06338_));
 sky130_fd_sc_hd__mux2_2 _12560_ (.A0(\core.cpuregs[8][14] ),
    .A1(\core.cpuregs[9][14] ),
    .S(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__mux2_2 _12561_ (.A0(\core.cpuregs[10][14] ),
    .A1(\core.cpuregs[11][14] ),
    .S(_06246_),
    .X(_06340_));
 sky130_fd_sc_hd__a21o_2 _12562_ (.A1(_06144_),
    .A2(_06340_),
    .B1(_06054_),
    .X(_06341_));
 sky130_fd_sc_hd__a21o_2 _12563_ (.A1(_06208_),
    .A2(_06339_),
    .B1(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__o211a_2 _12564_ (.A1(_06043_),
    .A2(_06337_),
    .B1(_06342_),
    .C1(_06058_),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_2 _12565_ (.A0(\core.cpuregs[4][14] ),
    .A1(\core.cpuregs[5][14] ),
    .S(_06062_),
    .X(_06344_));
 sky130_fd_sc_hd__and2_2 _12566_ (.A(_06149_),
    .B(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__mux2_2 _12567_ (.A0(\core.cpuregs[6][14] ),
    .A1(\core.cpuregs[7][14] ),
    .S(_06282_),
    .X(_06346_));
 sky130_fd_sc_hd__and2_2 _12568_ (.A(_06066_),
    .B(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__buf_1 _12569_ (.A(_02143_),
    .X(_06348_));
 sky130_fd_sc_hd__mux4_2 _12570_ (.A0(\core.cpuregs[0][14] ),
    .A1(\core.cpuregs[1][14] ),
    .A2(\core.cpuregs[2][14] ),
    .A3(\core.cpuregs[3][14] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06349_));
 sky130_fd_sc_hd__or2_2 _12571_ (.A(_06348_),
    .B(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__o311a_2 _12572_ (.A1(_06214_),
    .A2(_06345_),
    .A3(_06347_),
    .B1(_06070_),
    .C1(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__buf_1 _12573_ (.A(_06015_),
    .X(_06352_));
 sky130_fd_sc_hd__mux4_2 _12574_ (.A0(\core.cpuregs[16][14] ),
    .A1(\core.cpuregs[17][14] ),
    .A2(\core.cpuregs[18][14] ),
    .A3(\core.cpuregs[19][14] ),
    .S0(_06352_),
    .S1(_06158_),
    .X(_06353_));
 sky130_fd_sc_hd__nor2_2 _12575_ (.A(_06224_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__buf_1 _12576_ (.A(_02167_),
    .X(_06355_));
 sky130_fd_sc_hd__mux2_2 _12577_ (.A0(\core.cpuregs[20][14] ),
    .A1(\core.cpuregs[21][14] ),
    .S(_06161_),
    .X(_06356_));
 sky130_fd_sc_hd__mux2_2 _12578_ (.A0(\core.cpuregs[22][14] ),
    .A1(\core.cpuregs[23][14] ),
    .S(_06293_),
    .X(_06357_));
 sky130_fd_sc_hd__a21o_2 _12579_ (.A1(_06292_),
    .A2(_06357_),
    .B1(_06324_),
    .X(_06358_));
 sky130_fd_sc_hd__a21oi_2 _12580_ (.A1(_06355_),
    .A2(_06356_),
    .B1(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__mux2_2 _12581_ (.A0(\core.cpuregs[28][14] ),
    .A1(\core.cpuregs[29][14] ),
    .S(_06231_),
    .X(_06360_));
 sky130_fd_sc_hd__buf_1 _12582_ (.A(_06027_),
    .X(_06361_));
 sky130_fd_sc_hd__mux2_2 _12583_ (.A0(\core.cpuregs[30][14] ),
    .A1(\core.cpuregs[31][14] ),
    .S(_06233_),
    .X(_06362_));
 sky130_fd_sc_hd__a21o_2 _12584_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06197_),
    .X(_06363_));
 sky130_fd_sc_hd__a21oi_2 _12585_ (.A1(_06091_),
    .A2(_06360_),
    .B1(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__mux4_2 _12586_ (.A0(\core.cpuregs[24][14] ),
    .A1(\core.cpuregs[25][14] ),
    .A2(\core.cpuregs[26][14] ),
    .A3(\core.cpuregs[27][14] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06365_));
 sky130_fd_sc_hd__buf_1 _12587_ (.A(_02152_),
    .X(_06366_));
 sky130_fd_sc_hd__o21ai_2 _12588_ (.A1(_06099_),
    .A2(_06365_),
    .B1(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__o32a_2 _12589_ (.A1(_06223_),
    .A2(_06354_),
    .A3(_06359_),
    .B1(_06364_),
    .B2(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__nand2_2 _12590_ (.A(_06222_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__o311a_2 _12591_ (.A1(_06041_),
    .A2(_06343_),
    .A3(_06351_),
    .B1(_06369_),
    .C1(_06107_),
    .X(_06370_));
 sky130_fd_sc_hd__a21o_2 _12592_ (.A1(\core.decoded_imm[14] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06371_));
 sky130_fd_sc_hd__o22a_2 _12593_ (.A1(\core.pcpi_rs2[14] ),
    .A2(_06040_),
    .B1(_06370_),
    .B2(_06371_),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_2 _12594_ (.A0(\core.cpuregs[12][15] ),
    .A1(\core.cpuregs[13][15] ),
    .A2(\core.cpuregs[14][15] ),
    .A3(\core.cpuregs[15][15] ),
    .S0(_06045_),
    .S1(_06206_),
    .X(_06372_));
 sky130_fd_sc_hd__mux2_2 _12595_ (.A0(\core.cpuregs[8][15] ),
    .A1(\core.cpuregs[9][15] ),
    .S(_06338_),
    .X(_06373_));
 sky130_fd_sc_hd__mux2_2 _12596_ (.A0(\core.cpuregs[10][15] ),
    .A1(\core.cpuregs[11][15] ),
    .S(_06246_),
    .X(_06374_));
 sky130_fd_sc_hd__a21o_2 _12597_ (.A1(_06144_),
    .A2(_06374_),
    .B1(_06054_),
    .X(_06375_));
 sky130_fd_sc_hd__a21o_2 _12598_ (.A1(_06208_),
    .A2(_06373_),
    .B1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__o211a_2 _12599_ (.A1(_06043_),
    .A2(_06372_),
    .B1(_06376_),
    .C1(_06058_),
    .X(_06377_));
 sky130_fd_sc_hd__mux2_2 _12600_ (.A0(\core.cpuregs[4][15] ),
    .A1(\core.cpuregs[5][15] ),
    .S(_06062_),
    .X(_06378_));
 sky130_fd_sc_hd__and2_2 _12601_ (.A(_06149_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__mux2_2 _12602_ (.A0(\core.cpuregs[6][15] ),
    .A1(\core.cpuregs[7][15] ),
    .S(_06282_),
    .X(_06380_));
 sky130_fd_sc_hd__and2_2 _12603_ (.A(_06066_),
    .B(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__mux4_2 _12604_ (.A0(\core.cpuregs[0][15] ),
    .A1(\core.cpuregs[1][15] ),
    .A2(\core.cpuregs[2][15] ),
    .A3(\core.cpuregs[3][15] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06382_));
 sky130_fd_sc_hd__or2_2 _12605_ (.A(_06348_),
    .B(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__o311a_2 _12606_ (.A1(_06214_),
    .A2(_06379_),
    .A3(_06381_),
    .B1(_06070_),
    .C1(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__mux4_2 _12607_ (.A0(\core.cpuregs[16][15] ),
    .A1(\core.cpuregs[17][15] ),
    .A2(\core.cpuregs[18][15] ),
    .A3(\core.cpuregs[19][15] ),
    .S0(_06352_),
    .S1(_06158_),
    .X(_06385_));
 sky130_fd_sc_hd__nor2_2 _12608_ (.A(_06224_),
    .B(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__mux2_2 _12609_ (.A0(\core.cpuregs[20][15] ),
    .A1(\core.cpuregs[21][15] ),
    .S(_06161_),
    .X(_06387_));
 sky130_fd_sc_hd__mux2_2 _12610_ (.A0(\core.cpuregs[22][15] ),
    .A1(\core.cpuregs[23][15] ),
    .S(_06293_),
    .X(_06388_));
 sky130_fd_sc_hd__a21o_2 _12611_ (.A1(_06292_),
    .A2(_06388_),
    .B1(_06324_),
    .X(_06389_));
 sky130_fd_sc_hd__a21oi_2 _12612_ (.A1(_06355_),
    .A2(_06387_),
    .B1(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__mux2_2 _12613_ (.A0(\core.cpuregs[28][15] ),
    .A1(\core.cpuregs[29][15] ),
    .S(_06231_),
    .X(_06391_));
 sky130_fd_sc_hd__mux2_2 _12614_ (.A0(\core.cpuregs[30][15] ),
    .A1(\core.cpuregs[31][15] ),
    .S(_06233_),
    .X(_06392_));
 sky130_fd_sc_hd__a21o_2 _12615_ (.A1(_06361_),
    .A2(_06392_),
    .B1(_06197_),
    .X(_06393_));
 sky130_fd_sc_hd__a21oi_2 _12616_ (.A1(_06091_),
    .A2(_06391_),
    .B1(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__mux4_2 _12617_ (.A0(\core.cpuregs[24][15] ),
    .A1(\core.cpuregs[25][15] ),
    .A2(\core.cpuregs[26][15] ),
    .A3(\core.cpuregs[27][15] ),
    .S0(_06237_),
    .S1(_06101_),
    .X(_06395_));
 sky130_fd_sc_hd__o21ai_2 _12618_ (.A1(_06099_),
    .A2(_06395_),
    .B1(_06366_),
    .Y(_06396_));
 sky130_fd_sc_hd__o32a_2 _12619_ (.A1(_06223_),
    .A2(_06386_),
    .A3(_06390_),
    .B1(_06394_),
    .B2(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__nand2_2 _12620_ (.A(_06222_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__o311a_2 _12621_ (.A1(_06041_),
    .A2(_06377_),
    .A3(_06384_),
    .B1(_06398_),
    .C1(_06107_),
    .X(_06399_));
 sky130_fd_sc_hd__a21o_2 _12622_ (.A1(\core.decoded_imm[15] ),
    .A2(_06109_),
    .B1(_06111_),
    .X(_06400_));
 sky130_fd_sc_hd__o22a_2 _12623_ (.A1(\core.pcpi_rs2[15] ),
    .A2(_06040_),
    .B1(_06399_),
    .B2(_06400_),
    .X(_00619_));
 sky130_fd_sc_hd__buf_1 _12624_ (.A(_05987_),
    .X(_06401_));
 sky130_fd_sc_hd__buf_1 _12625_ (.A(_02127_),
    .X(_06402_));
 sky130_fd_sc_hd__buf_1 _12626_ (.A(_06042_),
    .X(_06403_));
 sky130_fd_sc_hd__buf_1 _12627_ (.A(_06044_),
    .X(_06404_));
 sky130_fd_sc_hd__mux4_2 _12628_ (.A0(\core.cpuregs[12][16] ),
    .A1(\core.cpuregs[13][16] ),
    .A2(\core.cpuregs[14][16] ),
    .A3(\core.cpuregs[15][16] ),
    .S0(_06404_),
    .S1(_06206_),
    .X(_06405_));
 sky130_fd_sc_hd__mux2_2 _12629_ (.A0(\core.cpuregs[8][16] ),
    .A1(\core.cpuregs[9][16] ),
    .S(_06338_),
    .X(_06406_));
 sky130_fd_sc_hd__mux2_2 _12630_ (.A0(\core.cpuregs[10][16] ),
    .A1(\core.cpuregs[11][16] ),
    .S(_06246_),
    .X(_06407_));
 sky130_fd_sc_hd__buf_1 _12631_ (.A(_02143_),
    .X(_06408_));
 sky130_fd_sc_hd__a21o_2 _12632_ (.A1(_06144_),
    .A2(_06407_),
    .B1(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__a21o_2 _12633_ (.A1(_06208_),
    .A2(_06406_),
    .B1(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__buf_1 _12634_ (.A(_06057_),
    .X(_06411_));
 sky130_fd_sc_hd__o211a_2 _12635_ (.A1(_06403_),
    .A2(_06405_),
    .B1(_06410_),
    .C1(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__buf_1 _12636_ (.A(_06018_),
    .X(_06413_));
 sky130_fd_sc_hd__mux2_2 _12637_ (.A0(\core.cpuregs[4][16] ),
    .A1(\core.cpuregs[5][16] ),
    .S(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__and2_2 _12638_ (.A(_06149_),
    .B(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__buf_1 _12639_ (.A(_06065_),
    .X(_06416_));
 sky130_fd_sc_hd__mux2_2 _12640_ (.A0(\core.cpuregs[6][16] ),
    .A1(\core.cpuregs[7][16] ),
    .S(_06282_),
    .X(_06417_));
 sky130_fd_sc_hd__and2_2 _12641_ (.A(_06416_),
    .B(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__buf_1 _12642_ (.A(_02129_),
    .X(_06419_));
 sky130_fd_sc_hd__mux4_2 _12643_ (.A0(\core.cpuregs[0][16] ),
    .A1(\core.cpuregs[1][16] ),
    .A2(\core.cpuregs[2][16] ),
    .A3(\core.cpuregs[3][16] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06420_));
 sky130_fd_sc_hd__or2_2 _12644_ (.A(_06348_),
    .B(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__o311a_2 _12645_ (.A1(_06214_),
    .A2(_06415_),
    .A3(_06418_),
    .B1(_06419_),
    .C1(_06421_),
    .X(_06422_));
 sky130_fd_sc_hd__mux4_2 _12646_ (.A0(\core.cpuregs[16][16] ),
    .A1(\core.cpuregs[17][16] ),
    .A2(\core.cpuregs[18][16] ),
    .A3(\core.cpuregs[19][16] ),
    .S0(_06352_),
    .S1(_06158_),
    .X(_06423_));
 sky130_fd_sc_hd__nor2_2 _12647_ (.A(_06224_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__mux2_2 _12648_ (.A0(\core.cpuregs[20][16] ),
    .A1(\core.cpuregs[21][16] ),
    .S(_06161_),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_2 _12649_ (.A0(\core.cpuregs[22][16] ),
    .A1(\core.cpuregs[23][16] ),
    .S(_06293_),
    .X(_06426_));
 sky130_fd_sc_hd__a21o_2 _12650_ (.A1(_06292_),
    .A2(_06426_),
    .B1(_06324_),
    .X(_06427_));
 sky130_fd_sc_hd__a21oi_2 _12651_ (.A1(_06355_),
    .A2(_06425_),
    .B1(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__buf_1 _12652_ (.A(_06024_),
    .X(_06429_));
 sky130_fd_sc_hd__mux2_2 _12653_ (.A0(\core.cpuregs[28][16] ),
    .A1(\core.cpuregs[29][16] ),
    .S(_06231_),
    .X(_06430_));
 sky130_fd_sc_hd__mux2_2 _12654_ (.A0(\core.cpuregs[30][16] ),
    .A1(\core.cpuregs[31][16] ),
    .S(_06233_),
    .X(_06431_));
 sky130_fd_sc_hd__a21o_2 _12655_ (.A1(_06361_),
    .A2(_06431_),
    .B1(_06197_),
    .X(_06432_));
 sky130_fd_sc_hd__a21oi_2 _12656_ (.A1(_06429_),
    .A2(_06430_),
    .B1(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__buf_1 _12657_ (.A(_06098_),
    .X(_06434_));
 sky130_fd_sc_hd__buf_1 _12658_ (.A(_06020_),
    .X(_06435_));
 sky130_fd_sc_hd__mux4_2 _12659_ (.A0(\core.cpuregs[24][16] ),
    .A1(\core.cpuregs[25][16] ),
    .A2(\core.cpuregs[26][16] ),
    .A3(\core.cpuregs[27][16] ),
    .S0(_06237_),
    .S1(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__o21ai_2 _12660_ (.A1(_06434_),
    .A2(_06436_),
    .B1(_06366_),
    .Y(_06437_));
 sky130_fd_sc_hd__o32a_2 _12661_ (.A1(_06223_),
    .A2(_06424_),
    .A3(_06428_),
    .B1(_06433_),
    .B2(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__nand2_2 _12662_ (.A(_06222_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__buf_1 _12663_ (.A(_05998_),
    .X(_06440_));
 sky130_fd_sc_hd__o311a_2 _12664_ (.A1(_06402_),
    .A2(_06412_),
    .A3(_06422_),
    .B1(_06439_),
    .C1(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_1 _12665_ (.A(_06037_),
    .X(_06442_));
 sky130_fd_sc_hd__buf_1 _12666_ (.A(_06110_),
    .X(_06443_));
 sky130_fd_sc_hd__a21o_2 _12667_ (.A1(\core.decoded_imm[16] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__o22a_2 _12668_ (.A1(\core.pcpi_rs2[16] ),
    .A2(_06401_),
    .B1(_06441_),
    .B2(_06444_),
    .X(_00620_));
 sky130_fd_sc_hd__mux4_2 _12669_ (.A0(\core.cpuregs[12][17] ),
    .A1(\core.cpuregs[13][17] ),
    .A2(\core.cpuregs[14][17] ),
    .A3(\core.cpuregs[15][17] ),
    .S0(_06404_),
    .S1(_06206_),
    .X(_06445_));
 sky130_fd_sc_hd__mux2_2 _12670_ (.A0(\core.cpuregs[8][17] ),
    .A1(\core.cpuregs[9][17] ),
    .S(_06338_),
    .X(_06446_));
 sky130_fd_sc_hd__mux2_2 _12671_ (.A0(\core.cpuregs[10][17] ),
    .A1(\core.cpuregs[11][17] ),
    .S(_06246_),
    .X(_06447_));
 sky130_fd_sc_hd__a21o_2 _12672_ (.A1(_06144_),
    .A2(_06447_),
    .B1(_06408_),
    .X(_06448_));
 sky130_fd_sc_hd__a21o_2 _12673_ (.A1(_06208_),
    .A2(_06446_),
    .B1(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__o211a_2 _12674_ (.A1(_06403_),
    .A2(_06445_),
    .B1(_06449_),
    .C1(_06411_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_2 _12675_ (.A0(\core.cpuregs[4][17] ),
    .A1(\core.cpuregs[5][17] ),
    .S(_06413_),
    .X(_06451_));
 sky130_fd_sc_hd__and2_2 _12676_ (.A(_06149_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__mux2_2 _12677_ (.A0(\core.cpuregs[6][17] ),
    .A1(\core.cpuregs[7][17] ),
    .S(_06282_),
    .X(_06453_));
 sky130_fd_sc_hd__and2_2 _12678_ (.A(_06416_),
    .B(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__mux4_2 _12679_ (.A0(\core.cpuregs[0][17] ),
    .A1(\core.cpuregs[1][17] ),
    .A2(\core.cpuregs[2][17] ),
    .A3(\core.cpuregs[3][17] ),
    .S0(_06154_),
    .S1(_06285_),
    .X(_06455_));
 sky130_fd_sc_hd__or2_2 _12680_ (.A(_06348_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__o311a_2 _12681_ (.A1(_06214_),
    .A2(_06452_),
    .A3(_06454_),
    .B1(_06419_),
    .C1(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__mux4_2 _12682_ (.A0(\core.cpuregs[16][17] ),
    .A1(\core.cpuregs[17][17] ),
    .A2(\core.cpuregs[18][17] ),
    .A3(\core.cpuregs[19][17] ),
    .S0(_06352_),
    .S1(_06158_),
    .X(_06458_));
 sky130_fd_sc_hd__nor2_2 _12683_ (.A(_06224_),
    .B(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__mux2_2 _12684_ (.A0(\core.cpuregs[20][17] ),
    .A1(\core.cpuregs[21][17] ),
    .S(_06161_),
    .X(_06460_));
 sky130_fd_sc_hd__mux2_2 _12685_ (.A0(\core.cpuregs[22][17] ),
    .A1(\core.cpuregs[23][17] ),
    .S(_06293_),
    .X(_06461_));
 sky130_fd_sc_hd__a21o_2 _12686_ (.A1(_06292_),
    .A2(_06461_),
    .B1(_06324_),
    .X(_06462_));
 sky130_fd_sc_hd__a21oi_2 _12687_ (.A1(_06355_),
    .A2(_06460_),
    .B1(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__mux2_2 _12688_ (.A0(\core.cpuregs[28][17] ),
    .A1(\core.cpuregs[29][17] ),
    .S(_06231_),
    .X(_06464_));
 sky130_fd_sc_hd__mux2_2 _12689_ (.A0(\core.cpuregs[30][17] ),
    .A1(\core.cpuregs[31][17] ),
    .S(_06233_),
    .X(_06465_));
 sky130_fd_sc_hd__a21o_2 _12690_ (.A1(_06361_),
    .A2(_06465_),
    .B1(_06197_),
    .X(_06466_));
 sky130_fd_sc_hd__a21oi_2 _12691_ (.A1(_06429_),
    .A2(_06464_),
    .B1(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__mux4_2 _12692_ (.A0(\core.cpuregs[24][17] ),
    .A1(\core.cpuregs[25][17] ),
    .A2(\core.cpuregs[26][17] ),
    .A3(\core.cpuregs[27][17] ),
    .S0(_06237_),
    .S1(_06435_),
    .X(_06468_));
 sky130_fd_sc_hd__o21ai_2 _12693_ (.A1(_06434_),
    .A2(_06468_),
    .B1(_06366_),
    .Y(_06469_));
 sky130_fd_sc_hd__o32a_2 _12694_ (.A1(_06223_),
    .A2(_06459_),
    .A3(_06463_),
    .B1(_06467_),
    .B2(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__nand2_2 _12695_ (.A(_06222_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__o311a_2 _12696_ (.A1(_06402_),
    .A2(_06450_),
    .A3(_06457_),
    .B1(_06471_),
    .C1(_06440_),
    .X(_06472_));
 sky130_fd_sc_hd__a21o_2 _12697_ (.A1(\core.decoded_imm[17] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06473_));
 sky130_fd_sc_hd__o22a_2 _12698_ (.A1(\core.pcpi_rs2[17] ),
    .A2(_06401_),
    .B1(_06472_),
    .B2(_06473_),
    .X(_00621_));
 sky130_fd_sc_hd__mux4_2 _12699_ (.A0(\core.cpuregs[12][18] ),
    .A1(\core.cpuregs[13][18] ),
    .A2(\core.cpuregs[14][18] ),
    .A3(\core.cpuregs[15][18] ),
    .S0(_06404_),
    .S1(_06206_),
    .X(_06474_));
 sky130_fd_sc_hd__mux2_2 _12700_ (.A0(\core.cpuregs[8][18] ),
    .A1(\core.cpuregs[9][18] ),
    .S(_06338_),
    .X(_06475_));
 sky130_fd_sc_hd__buf_1 _12701_ (.A(_06027_),
    .X(_06476_));
 sky130_fd_sc_hd__mux2_2 _12702_ (.A0(\core.cpuregs[10][18] ),
    .A1(\core.cpuregs[11][18] ),
    .S(_06246_),
    .X(_06477_));
 sky130_fd_sc_hd__a21o_2 _12703_ (.A1(_06476_),
    .A2(_06477_),
    .B1(_06408_),
    .X(_06478_));
 sky130_fd_sc_hd__a21o_2 _12704_ (.A1(_06208_),
    .A2(_06475_),
    .B1(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__o211a_2 _12705_ (.A1(_06403_),
    .A2(_06474_),
    .B1(_06479_),
    .C1(_06411_),
    .X(_06480_));
 sky130_fd_sc_hd__buf_1 _12706_ (.A(_02167_),
    .X(_06481_));
 sky130_fd_sc_hd__mux2_2 _12707_ (.A0(\core.cpuregs[4][18] ),
    .A1(\core.cpuregs[5][18] ),
    .S(_06413_),
    .X(_06482_));
 sky130_fd_sc_hd__and2_2 _12708_ (.A(_06481_),
    .B(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__mux2_2 _12709_ (.A0(\core.cpuregs[6][18] ),
    .A1(\core.cpuregs[7][18] ),
    .S(_06282_),
    .X(_06484_));
 sky130_fd_sc_hd__and2_2 _12710_ (.A(_06416_),
    .B(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__buf_1 _12711_ (.A(_06015_),
    .X(_06486_));
 sky130_fd_sc_hd__mux4_2 _12712_ (.A0(\core.cpuregs[0][18] ),
    .A1(\core.cpuregs[1][18] ),
    .A2(\core.cpuregs[2][18] ),
    .A3(\core.cpuregs[3][18] ),
    .S0(_06486_),
    .S1(_06285_),
    .X(_06487_));
 sky130_fd_sc_hd__or2_2 _12713_ (.A(_06348_),
    .B(_06487_),
    .X(_06488_));
 sky130_fd_sc_hd__o311a_2 _12714_ (.A1(_06214_),
    .A2(_06483_),
    .A3(_06485_),
    .B1(_06419_),
    .C1(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__buf_1 _12715_ (.A(_06020_),
    .X(_06490_));
 sky130_fd_sc_hd__mux4_2 _12716_ (.A0(\core.cpuregs[16][18] ),
    .A1(\core.cpuregs[17][18] ),
    .A2(\core.cpuregs[18][18] ),
    .A3(\core.cpuregs[19][18] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__nor2_2 _12717_ (.A(_06224_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__buf_1 _12718_ (.A(_06018_),
    .X(_06493_));
 sky130_fd_sc_hd__mux2_2 _12719_ (.A0(\core.cpuregs[20][18] ),
    .A1(\core.cpuregs[21][18] ),
    .S(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__mux2_2 _12720_ (.A0(\core.cpuregs[22][18] ),
    .A1(\core.cpuregs[23][18] ),
    .S(_06293_),
    .X(_06495_));
 sky130_fd_sc_hd__a21o_2 _12721_ (.A1(_06292_),
    .A2(_06495_),
    .B1(_06324_),
    .X(_06496_));
 sky130_fd_sc_hd__a21oi_2 _12722_ (.A1(_06355_),
    .A2(_06494_),
    .B1(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__mux2_2 _12723_ (.A0(\core.cpuregs[28][18] ),
    .A1(\core.cpuregs[29][18] ),
    .S(_06231_),
    .X(_06498_));
 sky130_fd_sc_hd__mux2_2 _12724_ (.A0(\core.cpuregs[30][18] ),
    .A1(\core.cpuregs[31][18] ),
    .S(_06233_),
    .X(_06499_));
 sky130_fd_sc_hd__a21o_2 _12725_ (.A1(_06361_),
    .A2(_06499_),
    .B1(_06197_),
    .X(_06500_));
 sky130_fd_sc_hd__a21oi_2 _12726_ (.A1(_06429_),
    .A2(_06498_),
    .B1(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__mux4_2 _12727_ (.A0(\core.cpuregs[24][18] ),
    .A1(\core.cpuregs[25][18] ),
    .A2(\core.cpuregs[26][18] ),
    .A3(\core.cpuregs[27][18] ),
    .S0(_06237_),
    .S1(_06435_),
    .X(_06502_));
 sky130_fd_sc_hd__o21ai_2 _12728_ (.A1(_06434_),
    .A2(_06502_),
    .B1(_06366_),
    .Y(_06503_));
 sky130_fd_sc_hd__o32a_2 _12729_ (.A1(_06223_),
    .A2(_06492_),
    .A3(_06497_),
    .B1(_06501_),
    .B2(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__nand2_2 _12730_ (.A(_06222_),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__o311a_2 _12731_ (.A1(_06402_),
    .A2(_06480_),
    .A3(_06489_),
    .B1(_06505_),
    .C1(_06440_),
    .X(_06506_));
 sky130_fd_sc_hd__a21o_2 _12732_ (.A1(\core.decoded_imm[18] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06507_));
 sky130_fd_sc_hd__o22a_2 _12733_ (.A1(\core.pcpi_rs2[18] ),
    .A2(_06401_),
    .B1(_06506_),
    .B2(_06507_),
    .X(_00622_));
 sky130_fd_sc_hd__mux4_2 _12734_ (.A0(\core.cpuregs[12][19] ),
    .A1(\core.cpuregs[13][19] ),
    .A2(\core.cpuregs[14][19] ),
    .A3(\core.cpuregs[15][19] ),
    .S0(_06404_),
    .S1(_06206_),
    .X(_06508_));
 sky130_fd_sc_hd__mux2_2 _12735_ (.A0(\core.cpuregs[8][19] ),
    .A1(\core.cpuregs[9][19] ),
    .S(_06338_),
    .X(_06509_));
 sky130_fd_sc_hd__mux2_2 _12736_ (.A0(\core.cpuregs[10][19] ),
    .A1(\core.cpuregs[11][19] ),
    .S(_06246_),
    .X(_06510_));
 sky130_fd_sc_hd__a21o_2 _12737_ (.A1(_06476_),
    .A2(_06510_),
    .B1(_06408_),
    .X(_06511_));
 sky130_fd_sc_hd__a21o_2 _12738_ (.A1(_06208_),
    .A2(_06509_),
    .B1(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__o211a_2 _12739_ (.A1(_06403_),
    .A2(_06508_),
    .B1(_06512_),
    .C1(_06411_),
    .X(_06513_));
 sky130_fd_sc_hd__mux2_2 _12740_ (.A0(\core.cpuregs[4][19] ),
    .A1(\core.cpuregs[5][19] ),
    .S(_06413_),
    .X(_06514_));
 sky130_fd_sc_hd__and2_2 _12741_ (.A(_06481_),
    .B(_06514_),
    .X(_06515_));
 sky130_fd_sc_hd__mux2_2 _12742_ (.A0(\core.cpuregs[6][19] ),
    .A1(\core.cpuregs[7][19] ),
    .S(_06282_),
    .X(_06516_));
 sky130_fd_sc_hd__and2_2 _12743_ (.A(_06416_),
    .B(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__mux4_2 _12744_ (.A0(\core.cpuregs[0][19] ),
    .A1(\core.cpuregs[1][19] ),
    .A2(\core.cpuregs[2][19] ),
    .A3(\core.cpuregs[3][19] ),
    .S0(_06486_),
    .S1(_06285_),
    .X(_06518_));
 sky130_fd_sc_hd__or2_2 _12745_ (.A(_06348_),
    .B(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__o311a_2 _12746_ (.A1(_06214_),
    .A2(_06515_),
    .A3(_06517_),
    .B1(_06419_),
    .C1(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__mux4_2 _12747_ (.A0(\core.cpuregs[16][19] ),
    .A1(\core.cpuregs[17][19] ),
    .A2(\core.cpuregs[18][19] ),
    .A3(\core.cpuregs[19][19] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06521_));
 sky130_fd_sc_hd__nor2_2 _12748_ (.A(_06224_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__mux2_2 _12749_ (.A0(\core.cpuregs[20][19] ),
    .A1(\core.cpuregs[21][19] ),
    .S(_06493_),
    .X(_06523_));
 sky130_fd_sc_hd__mux2_2 _12750_ (.A0(\core.cpuregs[22][19] ),
    .A1(\core.cpuregs[23][19] ),
    .S(_06293_),
    .X(_06524_));
 sky130_fd_sc_hd__a21o_2 _12751_ (.A1(_06292_),
    .A2(_06524_),
    .B1(_06324_),
    .X(_06525_));
 sky130_fd_sc_hd__a21oi_2 _12752_ (.A1(_06355_),
    .A2(_06523_),
    .B1(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__mux2_2 _12753_ (.A0(\core.cpuregs[28][19] ),
    .A1(\core.cpuregs[29][19] ),
    .S(_06231_),
    .X(_06527_));
 sky130_fd_sc_hd__mux2_2 _12754_ (.A0(\core.cpuregs[30][19] ),
    .A1(\core.cpuregs[31][19] ),
    .S(_06233_),
    .X(_06528_));
 sky130_fd_sc_hd__buf_1 _12755_ (.A(_02147_),
    .X(_06529_));
 sky130_fd_sc_hd__a21o_2 _12756_ (.A1(_06361_),
    .A2(_06528_),
    .B1(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__a21oi_2 _12757_ (.A1(_06429_),
    .A2(_06527_),
    .B1(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__mux4_2 _12758_ (.A0(\core.cpuregs[24][19] ),
    .A1(\core.cpuregs[25][19] ),
    .A2(\core.cpuregs[26][19] ),
    .A3(\core.cpuregs[27][19] ),
    .S0(_06237_),
    .S1(_06435_),
    .X(_06532_));
 sky130_fd_sc_hd__o21ai_2 _12759_ (.A1(_06434_),
    .A2(_06532_),
    .B1(_06366_),
    .Y(_06533_));
 sky130_fd_sc_hd__o32a_2 _12760_ (.A1(_06223_),
    .A2(_06522_),
    .A3(_06526_),
    .B1(_06531_),
    .B2(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__nand2_2 _12761_ (.A(_06222_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__o311a_2 _12762_ (.A1(_06402_),
    .A2(_06513_),
    .A3(_06520_),
    .B1(_06535_),
    .C1(_06440_),
    .X(_06536_));
 sky130_fd_sc_hd__a21o_2 _12763_ (.A1(\core.decoded_imm[19] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06537_));
 sky130_fd_sc_hd__o22a_2 _12764_ (.A1(\core.pcpi_rs2[19] ),
    .A2(_06401_),
    .B1(_06536_),
    .B2(_06537_),
    .X(_00623_));
 sky130_fd_sc_hd__buf_1 _12765_ (.A(_06027_),
    .X(_06538_));
 sky130_fd_sc_hd__mux4_2 _12766_ (.A0(\core.cpuregs[12][20] ),
    .A1(\core.cpuregs[13][20] ),
    .A2(\core.cpuregs[14][20] ),
    .A3(\core.cpuregs[15][20] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__buf_1 _12767_ (.A(_06024_),
    .X(_06540_));
 sky130_fd_sc_hd__mux2_2 _12768_ (.A0(\core.cpuregs[8][20] ),
    .A1(\core.cpuregs[9][20] ),
    .S(_06338_),
    .X(_06541_));
 sky130_fd_sc_hd__mux2_2 _12769_ (.A0(\core.cpuregs[10][20] ),
    .A1(\core.cpuregs[11][20] ),
    .S(_06246_),
    .X(_06542_));
 sky130_fd_sc_hd__a21o_2 _12770_ (.A1(_06476_),
    .A2(_06542_),
    .B1(_06408_),
    .X(_06543_));
 sky130_fd_sc_hd__a21o_2 _12771_ (.A1(_06540_),
    .A2(_06541_),
    .B1(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__o211a_2 _12772_ (.A1(_06403_),
    .A2(_06539_),
    .B1(_06544_),
    .C1(_06411_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_1 _12773_ (.A(_06042_),
    .X(_06546_));
 sky130_fd_sc_hd__mux2_2 _12774_ (.A0(\core.cpuregs[4][20] ),
    .A1(\core.cpuregs[5][20] ),
    .S(_06413_),
    .X(_06547_));
 sky130_fd_sc_hd__and2_2 _12775_ (.A(_06481_),
    .B(_06547_),
    .X(_06548_));
 sky130_fd_sc_hd__mux2_2 _12776_ (.A0(\core.cpuregs[6][20] ),
    .A1(\core.cpuregs[7][20] ),
    .S(_06282_),
    .X(_06549_));
 sky130_fd_sc_hd__and2_2 _12777_ (.A(_06416_),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__mux4_2 _12778_ (.A0(\core.cpuregs[0][20] ),
    .A1(\core.cpuregs[1][20] ),
    .A2(\core.cpuregs[2][20] ),
    .A3(\core.cpuregs[3][20] ),
    .S0(_06486_),
    .S1(_06285_),
    .X(_06551_));
 sky130_fd_sc_hd__or2_2 _12779_ (.A(_06348_),
    .B(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__o311a_2 _12780_ (.A1(_06546_),
    .A2(_06548_),
    .A3(_06550_),
    .B1(_06419_),
    .C1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__buf_1 _12781_ (.A(_02127_),
    .X(_06554_));
 sky130_fd_sc_hd__buf_1 _12782_ (.A(_02152_),
    .X(_06555_));
 sky130_fd_sc_hd__buf_1 _12783_ (.A(_06031_),
    .X(_06556_));
 sky130_fd_sc_hd__mux4_2 _12784_ (.A0(\core.cpuregs[16][20] ),
    .A1(\core.cpuregs[17][20] ),
    .A2(\core.cpuregs[18][20] ),
    .A3(\core.cpuregs[19][20] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06557_));
 sky130_fd_sc_hd__nor2_2 _12785_ (.A(_06556_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__mux2_2 _12786_ (.A0(\core.cpuregs[20][20] ),
    .A1(\core.cpuregs[21][20] ),
    .S(_06493_),
    .X(_06559_));
 sky130_fd_sc_hd__mux2_2 _12787_ (.A0(\core.cpuregs[22][20] ),
    .A1(\core.cpuregs[23][20] ),
    .S(_06293_),
    .X(_06560_));
 sky130_fd_sc_hd__a21o_2 _12788_ (.A1(_06292_),
    .A2(_06560_),
    .B1(_06324_),
    .X(_06561_));
 sky130_fd_sc_hd__a21oi_2 _12789_ (.A1(_06355_),
    .A2(_06559_),
    .B1(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__buf_1 _12790_ (.A(_06052_),
    .X(_06563_));
 sky130_fd_sc_hd__mux2_2 _12791_ (.A0(\core.cpuregs[28][20] ),
    .A1(\core.cpuregs[29][20] ),
    .S(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__buf_1 _12792_ (.A(_06000_),
    .X(_06565_));
 sky130_fd_sc_hd__mux2_2 _12793_ (.A0(\core.cpuregs[30][20] ),
    .A1(\core.cpuregs[31][20] ),
    .S(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__a21o_2 _12794_ (.A1(_06361_),
    .A2(_06566_),
    .B1(_06529_),
    .X(_06567_));
 sky130_fd_sc_hd__a21oi_2 _12795_ (.A1(_06429_),
    .A2(_06564_),
    .B1(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__buf_1 _12796_ (.A(_06015_),
    .X(_06569_));
 sky130_fd_sc_hd__mux4_2 _12797_ (.A0(\core.cpuregs[24][20] ),
    .A1(\core.cpuregs[25][20] ),
    .A2(\core.cpuregs[26][20] ),
    .A3(\core.cpuregs[27][20] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06570_));
 sky130_fd_sc_hd__o21ai_2 _12798_ (.A1(_06434_),
    .A2(_06570_),
    .B1(_06366_),
    .Y(_06571_));
 sky130_fd_sc_hd__o32a_2 _12799_ (.A1(_06555_),
    .A2(_06558_),
    .A3(_06562_),
    .B1(_06568_),
    .B2(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__nand2_2 _12800_ (.A(_06554_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__o311a_2 _12801_ (.A1(_06402_),
    .A2(_06545_),
    .A3(_06553_),
    .B1(_06573_),
    .C1(_06440_),
    .X(_06574_));
 sky130_fd_sc_hd__a21o_2 _12802_ (.A1(\core.decoded_imm[20] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06575_));
 sky130_fd_sc_hd__o22a_2 _12803_ (.A1(\core.pcpi_rs2[20] ),
    .A2(_06401_),
    .B1(_06574_),
    .B2(_06575_),
    .X(_00624_));
 sky130_fd_sc_hd__mux4_2 _12804_ (.A0(\core.cpuregs[12][21] ),
    .A1(\core.cpuregs[13][21] ),
    .A2(\core.cpuregs[14][21] ),
    .A3(\core.cpuregs[15][21] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06576_));
 sky130_fd_sc_hd__mux2_2 _12805_ (.A0(\core.cpuregs[8][21] ),
    .A1(\core.cpuregs[9][21] ),
    .S(_06338_),
    .X(_06577_));
 sky130_fd_sc_hd__buf_1 _12806_ (.A(_06000_),
    .X(_06578_));
 sky130_fd_sc_hd__mux2_2 _12807_ (.A0(\core.cpuregs[10][21] ),
    .A1(\core.cpuregs[11][21] ),
    .S(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__a21o_2 _12808_ (.A1(_06476_),
    .A2(_06579_),
    .B1(_06408_),
    .X(_06580_));
 sky130_fd_sc_hd__a21o_2 _12809_ (.A1(_06540_),
    .A2(_06577_),
    .B1(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__o211a_2 _12810_ (.A1(_06403_),
    .A2(_06576_),
    .B1(_06581_),
    .C1(_06411_),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_2 _12811_ (.A0(\core.cpuregs[4][21] ),
    .A1(\core.cpuregs[5][21] ),
    .S(_06413_),
    .X(_06583_));
 sky130_fd_sc_hd__and2_2 _12812_ (.A(_06481_),
    .B(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__mux2_2 _12813_ (.A0(\core.cpuregs[6][21] ),
    .A1(\core.cpuregs[7][21] ),
    .S(_06282_),
    .X(_06585_));
 sky130_fd_sc_hd__and2_2 _12814_ (.A(_06416_),
    .B(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__mux4_2 _12815_ (.A0(\core.cpuregs[0][21] ),
    .A1(\core.cpuregs[1][21] ),
    .A2(\core.cpuregs[2][21] ),
    .A3(\core.cpuregs[3][21] ),
    .S0(_06486_),
    .S1(_06285_),
    .X(_06587_));
 sky130_fd_sc_hd__or2_2 _12816_ (.A(_06348_),
    .B(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__o311a_2 _12817_ (.A1(_06546_),
    .A2(_06584_),
    .A3(_06586_),
    .B1(_06419_),
    .C1(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__mux4_2 _12818_ (.A0(\core.cpuregs[16][21] ),
    .A1(\core.cpuregs[17][21] ),
    .A2(\core.cpuregs[18][21] ),
    .A3(\core.cpuregs[19][21] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06590_));
 sky130_fd_sc_hd__nor2_2 _12819_ (.A(_06556_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__mux2_2 _12820_ (.A0(\core.cpuregs[20][21] ),
    .A1(\core.cpuregs[21][21] ),
    .S(_06493_),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_2 _12821_ (.A0(\core.cpuregs[22][21] ),
    .A1(\core.cpuregs[23][21] ),
    .S(_06293_),
    .X(_06593_));
 sky130_fd_sc_hd__a21o_2 _12822_ (.A1(_06292_),
    .A2(_06593_),
    .B1(_06324_),
    .X(_06594_));
 sky130_fd_sc_hd__a21oi_2 _12823_ (.A1(_06355_),
    .A2(_06592_),
    .B1(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__mux2_2 _12824_ (.A0(\core.cpuregs[28][21] ),
    .A1(\core.cpuregs[29][21] ),
    .S(_06563_),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_2 _12825_ (.A0(\core.cpuregs[30][21] ),
    .A1(\core.cpuregs[31][21] ),
    .S(_06565_),
    .X(_06597_));
 sky130_fd_sc_hd__a21o_2 _12826_ (.A1(_06361_),
    .A2(_06597_),
    .B1(_06529_),
    .X(_06598_));
 sky130_fd_sc_hd__a21oi_2 _12827_ (.A1(_06429_),
    .A2(_06596_),
    .B1(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__mux4_2 _12828_ (.A0(\core.cpuregs[24][21] ),
    .A1(\core.cpuregs[25][21] ),
    .A2(\core.cpuregs[26][21] ),
    .A3(\core.cpuregs[27][21] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06600_));
 sky130_fd_sc_hd__o21ai_2 _12829_ (.A1(_06434_),
    .A2(_06600_),
    .B1(_06366_),
    .Y(_06601_));
 sky130_fd_sc_hd__o32a_2 _12830_ (.A1(_06555_),
    .A2(_06591_),
    .A3(_06595_),
    .B1(_06599_),
    .B2(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__nand2_2 _12831_ (.A(_06554_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__o311a_2 _12832_ (.A1(_06402_),
    .A2(_06582_),
    .A3(_06589_),
    .B1(_06603_),
    .C1(_06440_),
    .X(_06604_));
 sky130_fd_sc_hd__a21o_2 _12833_ (.A1(\core.decoded_imm[21] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06605_));
 sky130_fd_sc_hd__o22a_2 _12834_ (.A1(\core.pcpi_rs2[21] ),
    .A2(_06401_),
    .B1(_06604_),
    .B2(_06605_),
    .X(_00625_));
 sky130_fd_sc_hd__mux4_2 _12835_ (.A0(\core.cpuregs[12][22] ),
    .A1(\core.cpuregs[13][22] ),
    .A2(\core.cpuregs[14][22] ),
    .A3(\core.cpuregs[15][22] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_2 _12836_ (.A0(\core.cpuregs[8][22] ),
    .A1(\core.cpuregs[9][22] ),
    .S(_06338_),
    .X(_06607_));
 sky130_fd_sc_hd__mux2_2 _12837_ (.A0(\core.cpuregs[10][22] ),
    .A1(\core.cpuregs[11][22] ),
    .S(_06578_),
    .X(_06608_));
 sky130_fd_sc_hd__a21o_2 _12838_ (.A1(_06476_),
    .A2(_06608_),
    .B1(_06408_),
    .X(_06609_));
 sky130_fd_sc_hd__a21o_2 _12839_ (.A1(_06540_),
    .A2(_06607_),
    .B1(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__o211a_2 _12840_ (.A1(_06403_),
    .A2(_06606_),
    .B1(_06610_),
    .C1(_06411_),
    .X(_06611_));
 sky130_fd_sc_hd__mux2_2 _12841_ (.A0(\core.cpuregs[4][22] ),
    .A1(\core.cpuregs[5][22] ),
    .S(_06413_),
    .X(_06612_));
 sky130_fd_sc_hd__and2_2 _12842_ (.A(_06481_),
    .B(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__buf_1 _12843_ (.A(_06018_),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_2 _12844_ (.A0(\core.cpuregs[6][22] ),
    .A1(\core.cpuregs[7][22] ),
    .S(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__and2_2 _12845_ (.A(_06416_),
    .B(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_1 _12846_ (.A(_02159_),
    .X(_06617_));
 sky130_fd_sc_hd__mux4_2 _12847_ (.A0(\core.cpuregs[0][22] ),
    .A1(\core.cpuregs[1][22] ),
    .A2(\core.cpuregs[2][22] ),
    .A3(\core.cpuregs[3][22] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__or2_2 _12848_ (.A(_06348_),
    .B(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__o311a_2 _12849_ (.A1(_06546_),
    .A2(_06613_),
    .A3(_06616_),
    .B1(_06419_),
    .C1(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__mux4_2 _12850_ (.A0(\core.cpuregs[16][22] ),
    .A1(\core.cpuregs[17][22] ),
    .A2(\core.cpuregs[18][22] ),
    .A3(\core.cpuregs[19][22] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06621_));
 sky130_fd_sc_hd__nor2_2 _12851_ (.A(_06556_),
    .B(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__mux2_2 _12852_ (.A0(\core.cpuregs[20][22] ),
    .A1(\core.cpuregs[21][22] ),
    .S(_06493_),
    .X(_06623_));
 sky130_fd_sc_hd__buf_1 _12853_ (.A(_06020_),
    .X(_06624_));
 sky130_fd_sc_hd__buf_1 _12854_ (.A(_06000_),
    .X(_06625_));
 sky130_fd_sc_hd__mux2_2 _12855_ (.A0(\core.cpuregs[22][22] ),
    .A1(\core.cpuregs[23][22] ),
    .S(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__a21o_2 _12856_ (.A1(_06624_),
    .A2(_06626_),
    .B1(_06324_),
    .X(_06627_));
 sky130_fd_sc_hd__a21oi_2 _12857_ (.A1(_06355_),
    .A2(_06623_),
    .B1(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__mux2_2 _12858_ (.A0(\core.cpuregs[28][22] ),
    .A1(\core.cpuregs[29][22] ),
    .S(_06563_),
    .X(_06629_));
 sky130_fd_sc_hd__mux2_2 _12859_ (.A0(\core.cpuregs[30][22] ),
    .A1(\core.cpuregs[31][22] ),
    .S(_06565_),
    .X(_06630_));
 sky130_fd_sc_hd__a21o_2 _12860_ (.A1(_06361_),
    .A2(_06630_),
    .B1(_06529_),
    .X(_06631_));
 sky130_fd_sc_hd__a21oi_2 _12861_ (.A1(_06429_),
    .A2(_06629_),
    .B1(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__mux4_2 _12862_ (.A0(\core.cpuregs[24][22] ),
    .A1(\core.cpuregs[25][22] ),
    .A2(\core.cpuregs[26][22] ),
    .A3(\core.cpuregs[27][22] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06633_));
 sky130_fd_sc_hd__o21ai_2 _12863_ (.A1(_06434_),
    .A2(_06633_),
    .B1(_06366_),
    .Y(_06634_));
 sky130_fd_sc_hd__o32a_2 _12864_ (.A1(_06555_),
    .A2(_06622_),
    .A3(_06628_),
    .B1(_06632_),
    .B2(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__nand2_2 _12865_ (.A(_06554_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__o311a_2 _12866_ (.A1(_06402_),
    .A2(_06611_),
    .A3(_06620_),
    .B1(_06636_),
    .C1(_06440_),
    .X(_06637_));
 sky130_fd_sc_hd__a21o_2 _12867_ (.A1(\core.decoded_imm[22] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06638_));
 sky130_fd_sc_hd__o22a_2 _12868_ (.A1(\core.pcpi_rs2[22] ),
    .A2(_06401_),
    .B1(_06637_),
    .B2(_06638_),
    .X(_00626_));
 sky130_fd_sc_hd__mux4_2 _12869_ (.A0(\core.cpuregs[12][23] ),
    .A1(\core.cpuregs[13][23] ),
    .A2(\core.cpuregs[14][23] ),
    .A3(\core.cpuregs[15][23] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06639_));
 sky130_fd_sc_hd__mux2_2 _12870_ (.A0(\core.cpuregs[8][23] ),
    .A1(\core.cpuregs[9][23] ),
    .S(_06338_),
    .X(_06640_));
 sky130_fd_sc_hd__mux2_2 _12871_ (.A0(\core.cpuregs[10][23] ),
    .A1(\core.cpuregs[11][23] ),
    .S(_06578_),
    .X(_06641_));
 sky130_fd_sc_hd__a21o_2 _12872_ (.A1(_06476_),
    .A2(_06641_),
    .B1(_06408_),
    .X(_06642_));
 sky130_fd_sc_hd__a21o_2 _12873_ (.A1(_06540_),
    .A2(_06640_),
    .B1(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__o211a_2 _12874_ (.A1(_06403_),
    .A2(_06639_),
    .B1(_06643_),
    .C1(_06411_),
    .X(_06644_));
 sky130_fd_sc_hd__mux2_2 _12875_ (.A0(\core.cpuregs[4][23] ),
    .A1(\core.cpuregs[5][23] ),
    .S(_06413_),
    .X(_06645_));
 sky130_fd_sc_hd__and2_2 _12876_ (.A(_06481_),
    .B(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__mux2_2 _12877_ (.A0(\core.cpuregs[6][23] ),
    .A1(\core.cpuregs[7][23] ),
    .S(_06614_),
    .X(_06647_));
 sky130_fd_sc_hd__and2_2 _12878_ (.A(_06416_),
    .B(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__mux4_2 _12879_ (.A0(\core.cpuregs[0][23] ),
    .A1(\core.cpuregs[1][23] ),
    .A2(\core.cpuregs[2][23] ),
    .A3(\core.cpuregs[3][23] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06649_));
 sky130_fd_sc_hd__or2_2 _12880_ (.A(_06348_),
    .B(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__o311a_2 _12881_ (.A1(_06546_),
    .A2(_06646_),
    .A3(_06648_),
    .B1(_06419_),
    .C1(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__mux4_2 _12882_ (.A0(\core.cpuregs[16][23] ),
    .A1(\core.cpuregs[17][23] ),
    .A2(\core.cpuregs[18][23] ),
    .A3(\core.cpuregs[19][23] ),
    .S0(_06352_),
    .S1(_06490_),
    .X(_06652_));
 sky130_fd_sc_hd__nor2_2 _12883_ (.A(_06556_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__mux2_2 _12884_ (.A0(\core.cpuregs[20][23] ),
    .A1(\core.cpuregs[21][23] ),
    .S(_06493_),
    .X(_06654_));
 sky130_fd_sc_hd__mux2_2 _12885_ (.A0(\core.cpuregs[22][23] ),
    .A1(\core.cpuregs[23][23] ),
    .S(_06625_),
    .X(_06655_));
 sky130_fd_sc_hd__a21o_2 _12886_ (.A1(_06624_),
    .A2(_06655_),
    .B1(_05999_),
    .X(_06656_));
 sky130_fd_sc_hd__a21oi_2 _12887_ (.A1(_06355_),
    .A2(_06654_),
    .B1(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__mux2_2 _12888_ (.A0(\core.cpuregs[28][23] ),
    .A1(\core.cpuregs[29][23] ),
    .S(_06563_),
    .X(_06658_));
 sky130_fd_sc_hd__mux2_2 _12889_ (.A0(\core.cpuregs[30][23] ),
    .A1(\core.cpuregs[31][23] ),
    .S(_06565_),
    .X(_06659_));
 sky130_fd_sc_hd__a21o_2 _12890_ (.A1(_06361_),
    .A2(_06659_),
    .B1(_06529_),
    .X(_06660_));
 sky130_fd_sc_hd__a21oi_2 _12891_ (.A1(_06429_),
    .A2(_06658_),
    .B1(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__mux4_2 _12892_ (.A0(\core.cpuregs[24][23] ),
    .A1(\core.cpuregs[25][23] ),
    .A2(\core.cpuregs[26][23] ),
    .A3(\core.cpuregs[27][23] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06662_));
 sky130_fd_sc_hd__o21ai_2 _12893_ (.A1(_06434_),
    .A2(_06662_),
    .B1(_06366_),
    .Y(_06663_));
 sky130_fd_sc_hd__o32a_2 _12894_ (.A1(_06555_),
    .A2(_06653_),
    .A3(_06657_),
    .B1(_06661_),
    .B2(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__nand2_2 _12895_ (.A(_06554_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__o311a_2 _12896_ (.A1(_06402_),
    .A2(_06644_),
    .A3(_06651_),
    .B1(_06665_),
    .C1(_06440_),
    .X(_06666_));
 sky130_fd_sc_hd__a21o_2 _12897_ (.A1(\core.decoded_imm[23] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06667_));
 sky130_fd_sc_hd__o22a_2 _12898_ (.A1(\core.pcpi_rs2[23] ),
    .A2(_06401_),
    .B1(_06666_),
    .B2(_06667_),
    .X(_00627_));
 sky130_fd_sc_hd__mux4_2 _12899_ (.A0(\core.cpuregs[12][24] ),
    .A1(\core.cpuregs[13][24] ),
    .A2(\core.cpuregs[14][24] ),
    .A3(\core.cpuregs[15][24] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06668_));
 sky130_fd_sc_hd__mux2_2 _12900_ (.A0(\core.cpuregs[8][24] ),
    .A1(\core.cpuregs[9][24] ),
    .S(_06084_),
    .X(_06669_));
 sky130_fd_sc_hd__mux2_2 _12901_ (.A0(\core.cpuregs[10][24] ),
    .A1(\core.cpuregs[11][24] ),
    .S(_06578_),
    .X(_06670_));
 sky130_fd_sc_hd__a21o_2 _12902_ (.A1(_06476_),
    .A2(_06670_),
    .B1(_06408_),
    .X(_06671_));
 sky130_fd_sc_hd__a21o_2 _12903_ (.A1(_06540_),
    .A2(_06669_),
    .B1(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__o211a_2 _12904_ (.A1(_06403_),
    .A2(_06668_),
    .B1(_06672_),
    .C1(_06411_),
    .X(_06673_));
 sky130_fd_sc_hd__mux2_2 _12905_ (.A0(\core.cpuregs[4][24] ),
    .A1(\core.cpuregs[5][24] ),
    .S(_06413_),
    .X(_06674_));
 sky130_fd_sc_hd__and2_2 _12906_ (.A(_06481_),
    .B(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__mux2_2 _12907_ (.A0(\core.cpuregs[6][24] ),
    .A1(\core.cpuregs[7][24] ),
    .S(_06614_),
    .X(_06676_));
 sky130_fd_sc_hd__and2_2 _12908_ (.A(_06416_),
    .B(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__mux4_2 _12909_ (.A0(\core.cpuregs[0][24] ),
    .A1(\core.cpuregs[1][24] ),
    .A2(\core.cpuregs[2][24] ),
    .A3(\core.cpuregs[3][24] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06678_));
 sky130_fd_sc_hd__or2_2 _12910_ (.A(_06098_),
    .B(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__o311a_2 _12911_ (.A1(_06546_),
    .A2(_06675_),
    .A3(_06677_),
    .B1(_06419_),
    .C1(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__mux4_2 _12912_ (.A0(\core.cpuregs[16][24] ),
    .A1(\core.cpuregs[17][24] ),
    .A2(\core.cpuregs[18][24] ),
    .A3(\core.cpuregs[19][24] ),
    .S0(_06072_),
    .S1(_06490_),
    .X(_06681_));
 sky130_fd_sc_hd__nor2_2 _12913_ (.A(_06556_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__mux2_2 _12914_ (.A0(\core.cpuregs[20][24] ),
    .A1(\core.cpuregs[21][24] ),
    .S(_06493_),
    .X(_06683_));
 sky130_fd_sc_hd__mux2_2 _12915_ (.A0(\core.cpuregs[22][24] ),
    .A1(\core.cpuregs[23][24] ),
    .S(_06625_),
    .X(_06684_));
 sky130_fd_sc_hd__a21o_2 _12916_ (.A1(_06624_),
    .A2(_06684_),
    .B1(_05999_),
    .X(_06685_));
 sky130_fd_sc_hd__a21oi_2 _12917_ (.A1(_06061_),
    .A2(_06683_),
    .B1(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__mux2_2 _12918_ (.A0(\core.cpuregs[28][24] ),
    .A1(\core.cpuregs[29][24] ),
    .S(_06563_),
    .X(_06687_));
 sky130_fd_sc_hd__mux2_2 _12919_ (.A0(\core.cpuregs[30][24] ),
    .A1(\core.cpuregs[31][24] ),
    .S(_06565_),
    .X(_06688_));
 sky130_fd_sc_hd__a21o_2 _12920_ (.A1(_06051_),
    .A2(_06688_),
    .B1(_06529_),
    .X(_06689_));
 sky130_fd_sc_hd__a21oi_2 _12921_ (.A1(_06429_),
    .A2(_06687_),
    .B1(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__mux4_2 _12922_ (.A0(\core.cpuregs[24][24] ),
    .A1(\core.cpuregs[25][24] ),
    .A2(\core.cpuregs[26][24] ),
    .A3(\core.cpuregs[27][24] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06691_));
 sky130_fd_sc_hd__o21ai_2 _12923_ (.A1(_06434_),
    .A2(_06691_),
    .B1(_06057_),
    .Y(_06692_));
 sky130_fd_sc_hd__o32a_2 _12924_ (.A1(_06555_),
    .A2(_06682_),
    .A3(_06686_),
    .B1(_06690_),
    .B2(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__nand2_2 _12925_ (.A(_06554_),
    .B(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__o311a_2 _12926_ (.A1(_06402_),
    .A2(_06673_),
    .A3(_06680_),
    .B1(_06694_),
    .C1(_06440_),
    .X(_06695_));
 sky130_fd_sc_hd__a21o_2 _12927_ (.A1(\core.decoded_imm[24] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06696_));
 sky130_fd_sc_hd__o22a_2 _12928_ (.A1(\core.pcpi_rs2[24] ),
    .A2(_06401_),
    .B1(_06695_),
    .B2(_06696_),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_2 _12929_ (.A0(\core.cpuregs[12][25] ),
    .A1(\core.cpuregs[13][25] ),
    .A2(\core.cpuregs[14][25] ),
    .A3(\core.cpuregs[15][25] ),
    .S0(_06404_),
    .S1(_06538_),
    .X(_06697_));
 sky130_fd_sc_hd__mux2_2 _12930_ (.A0(\core.cpuregs[8][25] ),
    .A1(\core.cpuregs[9][25] ),
    .S(_06084_),
    .X(_06698_));
 sky130_fd_sc_hd__mux2_2 _12931_ (.A0(\core.cpuregs[10][25] ),
    .A1(\core.cpuregs[11][25] ),
    .S(_06578_),
    .X(_06699_));
 sky130_fd_sc_hd__a21o_2 _12932_ (.A1(_06476_),
    .A2(_06699_),
    .B1(_06408_),
    .X(_06700_));
 sky130_fd_sc_hd__a21o_2 _12933_ (.A1(_06540_),
    .A2(_06698_),
    .B1(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__o211a_2 _12934_ (.A1(_06403_),
    .A2(_06697_),
    .B1(_06701_),
    .C1(_06411_),
    .X(_06702_));
 sky130_fd_sc_hd__mux2_2 _12935_ (.A0(\core.cpuregs[4][25] ),
    .A1(\core.cpuregs[5][25] ),
    .S(_06413_),
    .X(_06703_));
 sky130_fd_sc_hd__and2_2 _12936_ (.A(_06481_),
    .B(_06703_),
    .X(_06704_));
 sky130_fd_sc_hd__mux2_2 _12937_ (.A0(\core.cpuregs[6][25] ),
    .A1(\core.cpuregs[7][25] ),
    .S(_06614_),
    .X(_06705_));
 sky130_fd_sc_hd__and2_2 _12938_ (.A(_06416_),
    .B(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__mux4_2 _12939_ (.A0(\core.cpuregs[0][25] ),
    .A1(\core.cpuregs[1][25] ),
    .A2(\core.cpuregs[2][25] ),
    .A3(\core.cpuregs[3][25] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06707_));
 sky130_fd_sc_hd__or2_2 _12940_ (.A(_06098_),
    .B(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__o311a_2 _12941_ (.A1(_06546_),
    .A2(_06704_),
    .A3(_06706_),
    .B1(_06419_),
    .C1(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__mux4_2 _12942_ (.A0(\core.cpuregs[16][25] ),
    .A1(\core.cpuregs[17][25] ),
    .A2(\core.cpuregs[18][25] ),
    .A3(\core.cpuregs[19][25] ),
    .S0(_06072_),
    .S1(_06490_),
    .X(_06710_));
 sky130_fd_sc_hd__nor2_2 _12943_ (.A(_06556_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__mux2_2 _12944_ (.A0(\core.cpuregs[20][25] ),
    .A1(\core.cpuregs[21][25] ),
    .S(_06493_),
    .X(_06712_));
 sky130_fd_sc_hd__mux2_2 _12945_ (.A0(\core.cpuregs[22][25] ),
    .A1(\core.cpuregs[23][25] ),
    .S(_06625_),
    .X(_06713_));
 sky130_fd_sc_hd__a21o_2 _12946_ (.A1(_06624_),
    .A2(_06713_),
    .B1(_05999_),
    .X(_06714_));
 sky130_fd_sc_hd__a21oi_2 _12947_ (.A1(_06061_),
    .A2(_06712_),
    .B1(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__mux2_2 _12948_ (.A0(\core.cpuregs[28][25] ),
    .A1(\core.cpuregs[29][25] ),
    .S(_06563_),
    .X(_06716_));
 sky130_fd_sc_hd__mux2_2 _12949_ (.A0(\core.cpuregs[30][25] ),
    .A1(\core.cpuregs[31][25] ),
    .S(_06565_),
    .X(_06717_));
 sky130_fd_sc_hd__a21o_2 _12950_ (.A1(_06051_),
    .A2(_06717_),
    .B1(_06529_),
    .X(_06718_));
 sky130_fd_sc_hd__a21oi_2 _12951_ (.A1(_06429_),
    .A2(_06716_),
    .B1(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__mux4_2 _12952_ (.A0(\core.cpuregs[24][25] ),
    .A1(\core.cpuregs[25][25] ),
    .A2(\core.cpuregs[26][25] ),
    .A3(\core.cpuregs[27][25] ),
    .S0(_06569_),
    .S1(_06435_),
    .X(_06720_));
 sky130_fd_sc_hd__o21ai_2 _12953_ (.A1(_06434_),
    .A2(_06720_),
    .B1(_06057_),
    .Y(_06721_));
 sky130_fd_sc_hd__o32a_2 _12954_ (.A1(_06555_),
    .A2(_06711_),
    .A3(_06715_),
    .B1(_06719_),
    .B2(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__nand2_2 _12955_ (.A(_06554_),
    .B(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__o311a_2 _12956_ (.A1(_06402_),
    .A2(_06702_),
    .A3(_06709_),
    .B1(_06723_),
    .C1(_06440_),
    .X(_06724_));
 sky130_fd_sc_hd__a21o_2 _12957_ (.A1(\core.decoded_imm[25] ),
    .A2(_06442_),
    .B1(_06443_),
    .X(_06725_));
 sky130_fd_sc_hd__o22a_2 _12958_ (.A1(\core.pcpi_rs2[25] ),
    .A2(_06401_),
    .B1(_06724_),
    .B2(_06725_),
    .X(_00629_));
 sky130_fd_sc_hd__mux4_2 _12959_ (.A0(\core.cpuregs[12][26] ),
    .A1(\core.cpuregs[13][26] ),
    .A2(\core.cpuregs[14][26] ),
    .A3(\core.cpuregs[15][26] ),
    .S0(_06092_),
    .S1(_06538_),
    .X(_06726_));
 sky130_fd_sc_hd__mux2_2 _12960_ (.A0(\core.cpuregs[8][26] ),
    .A1(\core.cpuregs[9][26] ),
    .S(_06084_),
    .X(_06727_));
 sky130_fd_sc_hd__mux2_2 _12961_ (.A0(\core.cpuregs[10][26] ),
    .A1(\core.cpuregs[11][26] ),
    .S(_06578_),
    .X(_06728_));
 sky130_fd_sc_hd__a21o_2 _12962_ (.A1(_06476_),
    .A2(_06728_),
    .B1(_06031_),
    .X(_06729_));
 sky130_fd_sc_hd__a21o_2 _12963_ (.A1(_06540_),
    .A2(_06727_),
    .B1(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__o211a_2 _12964_ (.A1(_06060_),
    .A2(_06726_),
    .B1(_06730_),
    .C1(_06078_),
    .X(_06731_));
 sky130_fd_sc_hd__mux2_2 _12965_ (.A0(\core.cpuregs[4][26] ),
    .A1(\core.cpuregs[5][26] ),
    .S(_06100_),
    .X(_06732_));
 sky130_fd_sc_hd__and2_2 _12966_ (.A(_06481_),
    .B(_06732_),
    .X(_06733_));
 sky130_fd_sc_hd__mux2_2 _12967_ (.A0(\core.cpuregs[6][26] ),
    .A1(\core.cpuregs[7][26] ),
    .S(_06614_),
    .X(_06734_));
 sky130_fd_sc_hd__and2_2 _12968_ (.A(_06046_),
    .B(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__mux4_2 _12969_ (.A0(\core.cpuregs[0][26] ),
    .A1(\core.cpuregs[1][26] ),
    .A2(\core.cpuregs[2][26] ),
    .A3(\core.cpuregs[3][26] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06736_));
 sky130_fd_sc_hd__or2_2 _12970_ (.A(_06098_),
    .B(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__o311a_2 _12971_ (.A1(_06546_),
    .A2(_06733_),
    .A3(_06735_),
    .B1(_02129_),
    .C1(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__mux4_2 _12972_ (.A0(\core.cpuregs[16][26] ),
    .A1(\core.cpuregs[17][26] ),
    .A2(\core.cpuregs[18][26] ),
    .A3(\core.cpuregs[19][26] ),
    .S0(_06072_),
    .S1(_06490_),
    .X(_06739_));
 sky130_fd_sc_hd__nor2_2 _12973_ (.A(_06556_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__mux2_2 _12974_ (.A0(\core.cpuregs[20][26] ),
    .A1(\core.cpuregs[21][26] ),
    .S(_06493_),
    .X(_06741_));
 sky130_fd_sc_hd__mux2_2 _12975_ (.A0(\core.cpuregs[22][26] ),
    .A1(\core.cpuregs[23][26] ),
    .S(_06625_),
    .X(_06742_));
 sky130_fd_sc_hd__a21o_2 _12976_ (.A1(_06624_),
    .A2(_06742_),
    .B1(_05999_),
    .X(_06743_));
 sky130_fd_sc_hd__a21oi_2 _12977_ (.A1(_06061_),
    .A2(_06741_),
    .B1(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__mux2_2 _12978_ (.A0(\core.cpuregs[28][26] ),
    .A1(\core.cpuregs[29][26] ),
    .S(_06563_),
    .X(_06745_));
 sky130_fd_sc_hd__mux2_2 _12979_ (.A0(\core.cpuregs[30][26] ),
    .A1(\core.cpuregs[31][26] ),
    .S(_06565_),
    .X(_06746_));
 sky130_fd_sc_hd__a21o_2 _12980_ (.A1(_06051_),
    .A2(_06746_),
    .B1(_06529_),
    .X(_06747_));
 sky130_fd_sc_hd__a21oi_2 _12981_ (.A1(_06048_),
    .A2(_06745_),
    .B1(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__mux4_2 _12982_ (.A0(\core.cpuregs[24][26] ),
    .A1(\core.cpuregs[25][26] ),
    .A2(\core.cpuregs[26][26] ),
    .A3(\core.cpuregs[27][26] ),
    .S0(_06569_),
    .S1(_06065_),
    .X(_06749_));
 sky130_fd_sc_hd__o21ai_2 _12983_ (.A1(_06079_),
    .A2(_06749_),
    .B1(_06057_),
    .Y(_06750_));
 sky130_fd_sc_hd__o32a_2 _12984_ (.A1(_06555_),
    .A2(_06740_),
    .A3(_06744_),
    .B1(_06748_),
    .B2(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__nand2_2 _12985_ (.A(_06554_),
    .B(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__o311a_2 _12986_ (.A1(_06077_),
    .A2(_06731_),
    .A3(_06738_),
    .B1(_06752_),
    .C1(_05998_),
    .X(_06753_));
 sky130_fd_sc_hd__a21o_2 _12987_ (.A1(\core.decoded_imm[26] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06754_));
 sky130_fd_sc_hd__o22a_2 _12988_ (.A1(\core.pcpi_rs2[26] ),
    .A2(_05987_),
    .B1(_06753_),
    .B2(_06754_),
    .X(_00630_));
 sky130_fd_sc_hd__mux4_2 _12989_ (.A0(\core.cpuregs[12][27] ),
    .A1(\core.cpuregs[13][27] ),
    .A2(\core.cpuregs[14][27] ),
    .A3(\core.cpuregs[15][27] ),
    .S0(_06092_),
    .S1(_06538_),
    .X(_06755_));
 sky130_fd_sc_hd__mux2_2 _12990_ (.A0(\core.cpuregs[8][27] ),
    .A1(\core.cpuregs[9][27] ),
    .S(_06084_),
    .X(_06756_));
 sky130_fd_sc_hd__mux2_2 _12991_ (.A0(\core.cpuregs[10][27] ),
    .A1(\core.cpuregs[11][27] ),
    .S(_06578_),
    .X(_06757_));
 sky130_fd_sc_hd__a21o_2 _12992_ (.A1(_06476_),
    .A2(_06757_),
    .B1(_06031_),
    .X(_06758_));
 sky130_fd_sc_hd__a21o_2 _12993_ (.A1(_06540_),
    .A2(_06756_),
    .B1(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__o211a_2 _12994_ (.A1(_06060_),
    .A2(_06755_),
    .B1(_06759_),
    .C1(_06078_),
    .X(_06760_));
 sky130_fd_sc_hd__mux2_2 _12995_ (.A0(\core.cpuregs[4][27] ),
    .A1(\core.cpuregs[5][27] ),
    .S(_06100_),
    .X(_06761_));
 sky130_fd_sc_hd__and2_2 _12996_ (.A(_06481_),
    .B(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__mux2_2 _12997_ (.A0(\core.cpuregs[6][27] ),
    .A1(\core.cpuregs[7][27] ),
    .S(_06614_),
    .X(_06763_));
 sky130_fd_sc_hd__and2_2 _12998_ (.A(_06046_),
    .B(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__mux4_2 _12999_ (.A0(\core.cpuregs[0][27] ),
    .A1(\core.cpuregs[1][27] ),
    .A2(\core.cpuregs[2][27] ),
    .A3(\core.cpuregs[3][27] ),
    .S0(_06486_),
    .S1(_06617_),
    .X(_06765_));
 sky130_fd_sc_hd__or2_2 _13000_ (.A(_06098_),
    .B(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__o311a_2 _13001_ (.A1(_06546_),
    .A2(_06762_),
    .A3(_06764_),
    .B1(_02129_),
    .C1(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__mux4_2 _13002_ (.A0(\core.cpuregs[16][27] ),
    .A1(\core.cpuregs[17][27] ),
    .A2(\core.cpuregs[18][27] ),
    .A3(\core.cpuregs[19][27] ),
    .S0(_06072_),
    .S1(_06490_),
    .X(_06768_));
 sky130_fd_sc_hd__nor2_2 _13003_ (.A(_06556_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__mux2_2 _13004_ (.A0(\core.cpuregs[20][27] ),
    .A1(\core.cpuregs[21][27] ),
    .S(_06493_),
    .X(_06770_));
 sky130_fd_sc_hd__mux2_2 _13005_ (.A0(\core.cpuregs[22][27] ),
    .A1(\core.cpuregs[23][27] ),
    .S(_06625_),
    .X(_06771_));
 sky130_fd_sc_hd__a21o_2 _13006_ (.A1(_06624_),
    .A2(_06771_),
    .B1(_05999_),
    .X(_06772_));
 sky130_fd_sc_hd__a21oi_2 _13007_ (.A1(_06061_),
    .A2(_06770_),
    .B1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__mux2_2 _13008_ (.A0(\core.cpuregs[28][27] ),
    .A1(\core.cpuregs[29][27] ),
    .S(_06563_),
    .X(_06774_));
 sky130_fd_sc_hd__mux2_2 _13009_ (.A0(\core.cpuregs[30][27] ),
    .A1(\core.cpuregs[31][27] ),
    .S(_06565_),
    .X(_06775_));
 sky130_fd_sc_hd__a21o_2 _13010_ (.A1(_06051_),
    .A2(_06775_),
    .B1(_06529_),
    .X(_06776_));
 sky130_fd_sc_hd__a21oi_2 _13011_ (.A1(_06048_),
    .A2(_06774_),
    .B1(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__mux4_2 _13012_ (.A0(\core.cpuregs[24][27] ),
    .A1(\core.cpuregs[25][27] ),
    .A2(\core.cpuregs[26][27] ),
    .A3(\core.cpuregs[27][27] ),
    .S0(_06569_),
    .S1(_06065_),
    .X(_06778_));
 sky130_fd_sc_hd__o21ai_2 _13013_ (.A1(_06079_),
    .A2(_06778_),
    .B1(_06057_),
    .Y(_06779_));
 sky130_fd_sc_hd__o32a_2 _13014_ (.A1(_06555_),
    .A2(_06769_),
    .A3(_06773_),
    .B1(_06777_),
    .B2(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__nand2_2 _13015_ (.A(_06554_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__o311a_2 _13016_ (.A1(_06077_),
    .A2(_06760_),
    .A3(_06767_),
    .B1(_06781_),
    .C1(_05998_),
    .X(_06782_));
 sky130_fd_sc_hd__a21o_2 _13017_ (.A1(\core.decoded_imm[27] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06783_));
 sky130_fd_sc_hd__o22a_2 _13018_ (.A1(\core.pcpi_rs2[27] ),
    .A2(_05987_),
    .B1(_06782_),
    .B2(_06783_),
    .X(_00631_));
 sky130_fd_sc_hd__mux4_2 _13019_ (.A0(\core.cpuregs[12][28] ),
    .A1(\core.cpuregs[13][28] ),
    .A2(\core.cpuregs[14][28] ),
    .A3(\core.cpuregs[15][28] ),
    .S0(_06092_),
    .S1(_06538_),
    .X(_06784_));
 sky130_fd_sc_hd__mux2_2 _13020_ (.A0(\core.cpuregs[8][28] ),
    .A1(\core.cpuregs[9][28] ),
    .S(_06084_),
    .X(_06785_));
 sky130_fd_sc_hd__mux2_2 _13021_ (.A0(\core.cpuregs[10][28] ),
    .A1(\core.cpuregs[11][28] ),
    .S(_06578_),
    .X(_06786_));
 sky130_fd_sc_hd__a21o_2 _13022_ (.A1(_06086_),
    .A2(_06786_),
    .B1(_06031_),
    .X(_06787_));
 sky130_fd_sc_hd__a21o_2 _13023_ (.A1(_06540_),
    .A2(_06785_),
    .B1(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__o211a_2 _13024_ (.A1(_06060_),
    .A2(_06784_),
    .B1(_06788_),
    .C1(_06078_),
    .X(_06789_));
 sky130_fd_sc_hd__mux2_2 _13025_ (.A0(\core.cpuregs[4][28] ),
    .A1(\core.cpuregs[5][28] ),
    .S(_06100_),
    .X(_06790_));
 sky130_fd_sc_hd__and2_2 _13026_ (.A(_06024_),
    .B(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__mux2_2 _13027_ (.A0(\core.cpuregs[6][28] ),
    .A1(\core.cpuregs[7][28] ),
    .S(_06614_),
    .X(_06792_));
 sky130_fd_sc_hd__and2_2 _13028_ (.A(_06046_),
    .B(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__mux4_2 _13029_ (.A0(\core.cpuregs[0][28] ),
    .A1(\core.cpuregs[1][28] ),
    .A2(\core.cpuregs[2][28] ),
    .A3(\core.cpuregs[3][28] ),
    .S0(_06044_),
    .S1(_06617_),
    .X(_06794_));
 sky130_fd_sc_hd__or2_2 _13030_ (.A(_06098_),
    .B(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__o311a_2 _13031_ (.A1(_06546_),
    .A2(_06791_),
    .A3(_06793_),
    .B1(_02129_),
    .C1(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__mux4_2 _13032_ (.A0(\core.cpuregs[16][28] ),
    .A1(\core.cpuregs[17][28] ),
    .A2(\core.cpuregs[18][28] ),
    .A3(\core.cpuregs[19][28] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06797_));
 sky130_fd_sc_hd__nor2_2 _13033_ (.A(_06556_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__mux2_2 _13034_ (.A0(\core.cpuregs[20][28] ),
    .A1(\core.cpuregs[21][28] ),
    .S(_06067_),
    .X(_06799_));
 sky130_fd_sc_hd__mux2_2 _13035_ (.A0(\core.cpuregs[22][28] ),
    .A1(\core.cpuregs[23][28] ),
    .S(_06625_),
    .X(_06800_));
 sky130_fd_sc_hd__a21o_2 _13036_ (.A1(_06624_),
    .A2(_06800_),
    .B1(_05999_),
    .X(_06801_));
 sky130_fd_sc_hd__a21oi_2 _13037_ (.A1(_06061_),
    .A2(_06799_),
    .B1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__mux2_2 _13038_ (.A0(\core.cpuregs[28][28] ),
    .A1(\core.cpuregs[29][28] ),
    .S(_06563_),
    .X(_06803_));
 sky130_fd_sc_hd__mux2_2 _13039_ (.A0(\core.cpuregs[30][28] ),
    .A1(\core.cpuregs[31][28] ),
    .S(_06565_),
    .X(_06804_));
 sky130_fd_sc_hd__a21o_2 _13040_ (.A1(_06051_),
    .A2(_06804_),
    .B1(_06529_),
    .X(_06805_));
 sky130_fd_sc_hd__a21oi_2 _13041_ (.A1(_06048_),
    .A2(_06803_),
    .B1(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__mux4_2 _13042_ (.A0(\core.cpuregs[24][28] ),
    .A1(\core.cpuregs[25][28] ),
    .A2(\core.cpuregs[26][28] ),
    .A3(\core.cpuregs[27][28] ),
    .S0(_06569_),
    .S1(_06065_),
    .X(_06807_));
 sky130_fd_sc_hd__o21ai_2 _13043_ (.A1(_06079_),
    .A2(_06807_),
    .B1(_06057_),
    .Y(_06808_));
 sky130_fd_sc_hd__o32a_2 _13044_ (.A1(_06555_),
    .A2(_06798_),
    .A3(_06802_),
    .B1(_06806_),
    .B2(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__nand2_2 _13045_ (.A(_06554_),
    .B(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__o311a_2 _13046_ (.A1(_06077_),
    .A2(_06789_),
    .A3(_06796_),
    .B1(_06810_),
    .C1(_05998_),
    .X(_06811_));
 sky130_fd_sc_hd__a21o_2 _13047_ (.A1(\core.decoded_imm[28] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06812_));
 sky130_fd_sc_hd__o22a_2 _13048_ (.A1(\core.pcpi_rs2[28] ),
    .A2(_05987_),
    .B1(_06811_),
    .B2(_06812_),
    .X(_00632_));
 sky130_fd_sc_hd__mux4_2 _13049_ (.A0(\core.cpuregs[12][29] ),
    .A1(\core.cpuregs[13][29] ),
    .A2(\core.cpuregs[14][29] ),
    .A3(\core.cpuregs[15][29] ),
    .S0(_06092_),
    .S1(_06538_),
    .X(_06813_));
 sky130_fd_sc_hd__mux2_2 _13050_ (.A0(\core.cpuregs[8][29] ),
    .A1(\core.cpuregs[9][29] ),
    .S(_06084_),
    .X(_06814_));
 sky130_fd_sc_hd__mux2_2 _13051_ (.A0(\core.cpuregs[10][29] ),
    .A1(\core.cpuregs[11][29] ),
    .S(_06578_),
    .X(_06815_));
 sky130_fd_sc_hd__a21o_2 _13052_ (.A1(_06086_),
    .A2(_06815_),
    .B1(_06031_),
    .X(_06816_));
 sky130_fd_sc_hd__a21o_2 _13053_ (.A1(_06540_),
    .A2(_06814_),
    .B1(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__o211a_2 _13054_ (.A1(_06060_),
    .A2(_06813_),
    .B1(_06817_),
    .C1(_06078_),
    .X(_06818_));
 sky130_fd_sc_hd__mux2_2 _13055_ (.A0(\core.cpuregs[4][29] ),
    .A1(\core.cpuregs[5][29] ),
    .S(_06100_),
    .X(_06819_));
 sky130_fd_sc_hd__and2_2 _13056_ (.A(_06024_),
    .B(_06819_),
    .X(_06820_));
 sky130_fd_sc_hd__mux2_2 _13057_ (.A0(\core.cpuregs[6][29] ),
    .A1(\core.cpuregs[7][29] ),
    .S(_06614_),
    .X(_06821_));
 sky130_fd_sc_hd__and2_2 _13058_ (.A(_06046_),
    .B(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__mux4_2 _13059_ (.A0(\core.cpuregs[0][29] ),
    .A1(\core.cpuregs[1][29] ),
    .A2(\core.cpuregs[2][29] ),
    .A3(\core.cpuregs[3][29] ),
    .S0(_06044_),
    .S1(_06617_),
    .X(_06823_));
 sky130_fd_sc_hd__or2_2 _13060_ (.A(_06098_),
    .B(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__o311a_2 _13061_ (.A1(_06546_),
    .A2(_06820_),
    .A3(_06822_),
    .B1(_02129_),
    .C1(_06824_),
    .X(_06825_));
 sky130_fd_sc_hd__mux4_2 _13062_ (.A0(\core.cpuregs[16][29] ),
    .A1(\core.cpuregs[17][29] ),
    .A2(\core.cpuregs[18][29] ),
    .A3(\core.cpuregs[19][29] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06826_));
 sky130_fd_sc_hd__nor2_2 _13063_ (.A(_06556_),
    .B(_06826_),
    .Y(_06827_));
 sky130_fd_sc_hd__mux2_2 _13064_ (.A0(\core.cpuregs[20][29] ),
    .A1(\core.cpuregs[21][29] ),
    .S(_06067_),
    .X(_06828_));
 sky130_fd_sc_hd__mux2_2 _13065_ (.A0(\core.cpuregs[22][29] ),
    .A1(\core.cpuregs[23][29] ),
    .S(_06625_),
    .X(_06829_));
 sky130_fd_sc_hd__a21o_2 _13066_ (.A1(_06624_),
    .A2(_06829_),
    .B1(_05999_),
    .X(_06830_));
 sky130_fd_sc_hd__a21oi_2 _13067_ (.A1(_06061_),
    .A2(_06828_),
    .B1(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__mux2_2 _13068_ (.A0(\core.cpuregs[28][29] ),
    .A1(\core.cpuregs[29][29] ),
    .S(_06563_),
    .X(_06832_));
 sky130_fd_sc_hd__mux2_2 _13069_ (.A0(\core.cpuregs[30][29] ),
    .A1(\core.cpuregs[31][29] ),
    .S(_06565_),
    .X(_06833_));
 sky130_fd_sc_hd__a21o_2 _13070_ (.A1(_06051_),
    .A2(_06833_),
    .B1(_06088_),
    .X(_06834_));
 sky130_fd_sc_hd__a21oi_2 _13071_ (.A1(_06048_),
    .A2(_06832_),
    .B1(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__mux4_2 _13072_ (.A0(\core.cpuregs[24][29] ),
    .A1(\core.cpuregs[25][29] ),
    .A2(\core.cpuregs[26][29] ),
    .A3(\core.cpuregs[27][29] ),
    .S0(_06569_),
    .S1(_06065_),
    .X(_06836_));
 sky130_fd_sc_hd__o21ai_2 _13073_ (.A1(_06079_),
    .A2(_06836_),
    .B1(_06057_),
    .Y(_06837_));
 sky130_fd_sc_hd__o32a_2 _13074_ (.A1(_06555_),
    .A2(_06827_),
    .A3(_06831_),
    .B1(_06835_),
    .B2(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__nand2_2 _13075_ (.A(_06554_),
    .B(_06838_),
    .Y(_06839_));
 sky130_fd_sc_hd__o311a_2 _13076_ (.A1(_06077_),
    .A2(_06818_),
    .A3(_06825_),
    .B1(_06839_),
    .C1(_05998_),
    .X(_06840_));
 sky130_fd_sc_hd__a21o_2 _13077_ (.A1(\core.decoded_imm[29] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06841_));
 sky130_fd_sc_hd__o22a_2 _13078_ (.A1(\core.pcpi_rs2[29] ),
    .A2(_05987_),
    .B1(_06840_),
    .B2(_06841_),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_2 _13079_ (.A0(\core.cpuregs[12][30] ),
    .A1(\core.cpuregs[13][30] ),
    .A2(\core.cpuregs[14][30] ),
    .A3(\core.cpuregs[15][30] ),
    .S0(_06092_),
    .S1(_06094_),
    .X(_06842_));
 sky130_fd_sc_hd__mux2_2 _13080_ (.A0(\core.cpuregs[8][30] ),
    .A1(\core.cpuregs[9][30] ),
    .S(_06084_),
    .X(_06843_));
 sky130_fd_sc_hd__mux2_2 _13081_ (.A0(\core.cpuregs[10][30] ),
    .A1(\core.cpuregs[11][30] ),
    .S(_06578_),
    .X(_06844_));
 sky130_fd_sc_hd__a21o_2 _13082_ (.A1(_06086_),
    .A2(_06844_),
    .B1(_06031_),
    .X(_06845_));
 sky130_fd_sc_hd__a21o_2 _13083_ (.A1(_06083_),
    .A2(_06843_),
    .B1(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__o211a_2 _13084_ (.A1(_06060_),
    .A2(_06842_),
    .B1(_06846_),
    .C1(_06078_),
    .X(_06847_));
 sky130_fd_sc_hd__mux2_2 _13085_ (.A0(\core.cpuregs[4][30] ),
    .A1(\core.cpuregs[5][30] ),
    .S(_06100_),
    .X(_06848_));
 sky130_fd_sc_hd__and2_2 _13086_ (.A(_06024_),
    .B(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__mux2_2 _13087_ (.A0(\core.cpuregs[6][30] ),
    .A1(\core.cpuregs[7][30] ),
    .S(_06614_),
    .X(_06850_));
 sky130_fd_sc_hd__and2_2 _13088_ (.A(_06046_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__mux4_2 _13089_ (.A0(\core.cpuregs[0][30] ),
    .A1(\core.cpuregs[1][30] ),
    .A2(\core.cpuregs[2][30] ),
    .A3(\core.cpuregs[3][30] ),
    .S0(_06044_),
    .S1(_06617_),
    .X(_06852_));
 sky130_fd_sc_hd__or2_2 _13090_ (.A(_06098_),
    .B(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__o311a_2 _13091_ (.A1(_06042_),
    .A2(_06849_),
    .A3(_06851_),
    .B1(_02129_),
    .C1(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__mux4_2 _13092_ (.A0(\core.cpuregs[16][30] ),
    .A1(\core.cpuregs[17][30] ),
    .A2(\core.cpuregs[18][30] ),
    .A3(\core.cpuregs[19][30] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06855_));
 sky130_fd_sc_hd__nor2_2 _13093_ (.A(_06071_),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__mux2_2 _13094_ (.A0(\core.cpuregs[20][30] ),
    .A1(\core.cpuregs[21][30] ),
    .S(_06067_),
    .X(_06857_));
 sky130_fd_sc_hd__mux2_2 _13095_ (.A0(\core.cpuregs[22][30] ),
    .A1(\core.cpuregs[23][30] ),
    .S(_06625_),
    .X(_06858_));
 sky130_fd_sc_hd__a21o_2 _13096_ (.A1(_06624_),
    .A2(_06858_),
    .B1(_05999_),
    .X(_06859_));
 sky130_fd_sc_hd__a21oi_2 _13097_ (.A1(_06061_),
    .A2(_06857_),
    .B1(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__mux2_2 _13098_ (.A0(\core.cpuregs[28][30] ),
    .A1(\core.cpuregs[29][30] ),
    .S(_06049_),
    .X(_06861_));
 sky130_fd_sc_hd__mux2_2 _13099_ (.A0(\core.cpuregs[30][30] ),
    .A1(\core.cpuregs[31][30] ),
    .S(_06052_),
    .X(_06862_));
 sky130_fd_sc_hd__a21o_2 _13100_ (.A1(_06051_),
    .A2(_06862_),
    .B1(_06088_),
    .X(_06863_));
 sky130_fd_sc_hd__a21oi_2 _13101_ (.A1(_06048_),
    .A2(_06861_),
    .B1(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__mux4_2 _13102_ (.A0(\core.cpuregs[24][30] ),
    .A1(\core.cpuregs[25][30] ),
    .A2(\core.cpuregs[26][30] ),
    .A3(\core.cpuregs[27][30] ),
    .S0(_06080_),
    .S1(_06065_),
    .X(_06865_));
 sky130_fd_sc_hd__o21ai_2 _13103_ (.A1(_06079_),
    .A2(_06865_),
    .B1(_06057_),
    .Y(_06866_));
 sky130_fd_sc_hd__o32a_2 _13104_ (.A1(_06103_),
    .A2(_06856_),
    .A3(_06860_),
    .B1(_06864_),
    .B2(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__nand2_2 _13105_ (.A(_02127_),
    .B(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__o311a_2 _13106_ (.A1(_06077_),
    .A2(_06847_),
    .A3(_06854_),
    .B1(_06868_),
    .C1(_05998_),
    .X(_06869_));
 sky130_fd_sc_hd__a21o_2 _13107_ (.A1(\core.decoded_imm[30] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06870_));
 sky130_fd_sc_hd__o22a_2 _13108_ (.A1(\core.pcpi_rs2[30] ),
    .A2(_05987_),
    .B1(_06869_),
    .B2(_06870_),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_2 _13109_ (.A0(\core.cpuregs[12][31] ),
    .A1(\core.cpuregs[13][31] ),
    .A2(\core.cpuregs[14][31] ),
    .A3(\core.cpuregs[15][31] ),
    .S0(_06092_),
    .S1(_06094_),
    .X(_06871_));
 sky130_fd_sc_hd__mux2_2 _13110_ (.A0(\core.cpuregs[8][31] ),
    .A1(\core.cpuregs[9][31] ),
    .S(_06084_),
    .X(_06872_));
 sky130_fd_sc_hd__mux2_2 _13111_ (.A0(\core.cpuregs[10][31] ),
    .A1(\core.cpuregs[11][31] ),
    .S(_06025_),
    .X(_06873_));
 sky130_fd_sc_hd__a21o_2 _13112_ (.A1(_06086_),
    .A2(_06873_),
    .B1(_06031_),
    .X(_06874_));
 sky130_fd_sc_hd__a21o_2 _13113_ (.A1(_06083_),
    .A2(_06872_),
    .B1(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__o211a_2 _13114_ (.A1(_06060_),
    .A2(_06871_),
    .B1(_06875_),
    .C1(_06078_),
    .X(_06876_));
 sky130_fd_sc_hd__mux2_2 _13115_ (.A0(\core.cpuregs[4][31] ),
    .A1(\core.cpuregs[5][31] ),
    .S(_06100_),
    .X(_06877_));
 sky130_fd_sc_hd__and2_2 _13116_ (.A(_06024_),
    .B(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__mux2_2 _13117_ (.A0(\core.cpuregs[6][31] ),
    .A1(\core.cpuregs[7][31] ),
    .S(_06614_),
    .X(_06879_));
 sky130_fd_sc_hd__and2_2 _13118_ (.A(_06046_),
    .B(_06879_),
    .X(_06880_));
 sky130_fd_sc_hd__mux4_2 _13119_ (.A0(\core.cpuregs[0][31] ),
    .A1(\core.cpuregs[1][31] ),
    .A2(\core.cpuregs[2][31] ),
    .A3(\core.cpuregs[3][31] ),
    .S0(_06044_),
    .S1(_06617_),
    .X(_06881_));
 sky130_fd_sc_hd__or2_2 _13120_ (.A(_06098_),
    .B(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__o311a_2 _13121_ (.A1(_06042_),
    .A2(_06878_),
    .A3(_06880_),
    .B1(_02129_),
    .C1(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__mux4_2 _13122_ (.A0(\core.cpuregs[16][31] ),
    .A1(\core.cpuregs[17][31] ),
    .A2(\core.cpuregs[18][31] ),
    .A3(\core.cpuregs[19][31] ),
    .S0(_06072_),
    .S1(_06073_),
    .X(_06884_));
 sky130_fd_sc_hd__nor2_2 _13123_ (.A(_06071_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__mux2_2 _13124_ (.A0(\core.cpuregs[20][31] ),
    .A1(\core.cpuregs[21][31] ),
    .S(_06067_),
    .X(_06886_));
 sky130_fd_sc_hd__mux2_2 _13125_ (.A0(\core.cpuregs[22][31] ),
    .A1(\core.cpuregs[23][31] ),
    .S(_06625_),
    .X(_06887_));
 sky130_fd_sc_hd__a21o_2 _13126_ (.A1(_06624_),
    .A2(_06887_),
    .B1(_05999_),
    .X(_06888_));
 sky130_fd_sc_hd__a21oi_2 _13127_ (.A1(_06061_),
    .A2(_06886_),
    .B1(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__mux2_2 _13128_ (.A0(\core.cpuregs[28][31] ),
    .A1(\core.cpuregs[29][31] ),
    .S(_06049_),
    .X(_06890_));
 sky130_fd_sc_hd__mux2_2 _13129_ (.A0(\core.cpuregs[30][31] ),
    .A1(\core.cpuregs[31][31] ),
    .S(_06052_),
    .X(_06891_));
 sky130_fd_sc_hd__a21o_2 _13130_ (.A1(_06051_),
    .A2(_06891_),
    .B1(_06088_),
    .X(_06892_));
 sky130_fd_sc_hd__a21oi_2 _13131_ (.A1(_06048_),
    .A2(_06890_),
    .B1(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__mux4_2 _13132_ (.A0(\core.cpuregs[24][31] ),
    .A1(\core.cpuregs[25][31] ),
    .A2(\core.cpuregs[26][31] ),
    .A3(\core.cpuregs[27][31] ),
    .S0(_06080_),
    .S1(_06065_),
    .X(_06894_));
 sky130_fd_sc_hd__o21ai_2 _13133_ (.A1(_06079_),
    .A2(_06894_),
    .B1(_06057_),
    .Y(_06895_));
 sky130_fd_sc_hd__o32a_2 _13134_ (.A1(_06103_),
    .A2(_06885_),
    .A3(_06889_),
    .B1(_06893_),
    .B2(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__nand2_2 _13135_ (.A(_02127_),
    .B(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__o311a_2 _13136_ (.A1(_06077_),
    .A2(_06876_),
    .A3(_06883_),
    .B1(_06897_),
    .C1(_05998_),
    .X(_06898_));
 sky130_fd_sc_hd__a21o_2 _13137_ (.A1(\core.decoded_imm[31] ),
    .A2(_06037_),
    .B1(_06110_),
    .X(_06899_));
 sky130_fd_sc_hd__o22a_2 _13138_ (.A1(\core.pcpi_rs2[31] ),
    .A2(_05987_),
    .B1(_06898_),
    .B2(_06899_),
    .X(_00635_));
 sky130_fd_sc_hd__and2_2 _13139_ (.A(_05877_),
    .B(_05953_),
    .X(_06900_));
 sky130_fd_sc_hd__a22o_2 _13140_ (.A1(\core.instr_bge ),
    .A2(_05932_),
    .B1(_06900_),
    .B2(_02236_),
    .X(_06901_));
 sky130_fd_sc_hd__and2_2 _13141_ (.A(_05928_),
    .B(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__buf_1 _13142_ (.A(_06902_),
    .X(_00636_));
 sky130_fd_sc_hd__nor2_2 _13143_ (.A(_02117_),
    .B(_05830_),
    .Y(_06903_));
 sky130_fd_sc_hd__a22o_2 _13144_ (.A1(\core.instr_bltu ),
    .A2(_05932_),
    .B1(_05933_),
    .B2(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__and2_2 _13145_ (.A(_05928_),
    .B(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__buf_1 _13146_ (.A(_06905_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_2 _13147_ (.A0(\core.mem_rdata_q[12] ),
    .A1(mem_rdata[12]),
    .S(_03176_),
    .X(_06906_));
 sky130_fd_sc_hd__buf_1 _13148_ (.A(_06906_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_2 _13149_ (.A0(\core.mem_rdata_q[13] ),
    .A1(mem_rdata[13]),
    .S(_03176_),
    .X(_06907_));
 sky130_fd_sc_hd__buf_1 _13150_ (.A(_06907_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_2 _13151_ (.A0(\core.mem_rdata_q[14] ),
    .A1(mem_rdata[14]),
    .S(_03176_),
    .X(_06908_));
 sky130_fd_sc_hd__buf_1 _13152_ (.A(_06908_),
    .X(_01357_));
 sky130_fd_sc_hd__nor3_2 _13153_ (.A(_01355_),
    .B(_01356_),
    .C(_01357_),
    .Y(_06909_));
 sky130_fd_sc_hd__a32o_2 _13154_ (.A1(_05816_),
    .A2(_05874_),
    .A3(_06909_),
    .B1(_05803_),
    .B2(\core.instr_jalr ),
    .X(_00638_));
 sky130_fd_sc_hd__a22o_2 _13155_ (.A1(\core.instr_lb ),
    .A2(_05921_),
    .B1(_05881_),
    .B2(_02091_),
    .X(_00639_));
 sky130_fd_sc_hd__nor2_2 _13156_ (.A(_05285_),
    .B(_05766_),
    .Y(_06910_));
 sky130_fd_sc_hd__buf_1 _13157_ (.A(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__mux2_2 _13158_ (.A0(\core.cpuregs[20][0] ),
    .A1(_05284_),
    .S(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__buf_1 _13159_ (.A(_06912_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_2 _13160_ (.A0(\core.cpuregs[20][1] ),
    .A1(_05292_),
    .S(_06911_),
    .X(_06913_));
 sky130_fd_sc_hd__buf_1 _13161_ (.A(_06913_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_2 _13162_ (.A0(\core.cpuregs[20][2] ),
    .A1(_05297_),
    .S(_06911_),
    .X(_06914_));
 sky130_fd_sc_hd__buf_1 _13163_ (.A(_06914_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_2 _13164_ (.A0(\core.cpuregs[20][3] ),
    .A1(_05304_),
    .S(_06911_),
    .X(_06915_));
 sky130_fd_sc_hd__buf_1 _13165_ (.A(_06915_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_2 _13166_ (.A0(\core.cpuregs[20][4] ),
    .A1(_05310_),
    .S(_06911_),
    .X(_06916_));
 sky130_fd_sc_hd__buf_1 _13167_ (.A(_06916_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_2 _13168_ (.A0(\core.cpuregs[20][5] ),
    .A1(_05315_),
    .S(_06911_),
    .X(_06917_));
 sky130_fd_sc_hd__buf_1 _13169_ (.A(_06917_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_2 _13170_ (.A0(\core.cpuregs[20][6] ),
    .A1(_05320_),
    .S(_06911_),
    .X(_06918_));
 sky130_fd_sc_hd__buf_1 _13171_ (.A(_06918_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_2 _13172_ (.A0(\core.cpuregs[20][7] ),
    .A1(_05326_),
    .S(_06911_),
    .X(_06919_));
 sky130_fd_sc_hd__buf_1 _13173_ (.A(_06919_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_2 _13174_ (.A0(\core.cpuregs[20][8] ),
    .A1(_05332_),
    .S(_06911_),
    .X(_06920_));
 sky130_fd_sc_hd__buf_1 _13175_ (.A(_06920_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_2 _13176_ (.A0(\core.cpuregs[20][9] ),
    .A1(_05337_),
    .S(_06911_),
    .X(_06921_));
 sky130_fd_sc_hd__buf_1 _13177_ (.A(_06921_),
    .X(_00649_));
 sky130_fd_sc_hd__buf_1 _13178_ (.A(_06910_),
    .X(_06922_));
 sky130_fd_sc_hd__mux2_2 _13179_ (.A0(\core.cpuregs[20][10] ),
    .A1(_05343_),
    .S(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__buf_1 _13180_ (.A(_06923_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_2 _13181_ (.A0(\core.cpuregs[20][11] ),
    .A1(_05349_),
    .S(_06922_),
    .X(_06924_));
 sky130_fd_sc_hd__buf_1 _13182_ (.A(_06924_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_2 _13183_ (.A0(\core.cpuregs[20][12] ),
    .A1(_05355_),
    .S(_06922_),
    .X(_06925_));
 sky130_fd_sc_hd__buf_1 _13184_ (.A(_06925_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_2 _13185_ (.A0(\core.cpuregs[20][13] ),
    .A1(_05360_),
    .S(_06922_),
    .X(_06926_));
 sky130_fd_sc_hd__buf_1 _13186_ (.A(_06926_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_2 _13187_ (.A0(\core.cpuregs[20][14] ),
    .A1(_05367_),
    .S(_06922_),
    .X(_06927_));
 sky130_fd_sc_hd__buf_1 _13188_ (.A(_06927_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_2 _13189_ (.A0(\core.cpuregs[20][15] ),
    .A1(_05372_),
    .S(_06922_),
    .X(_06928_));
 sky130_fd_sc_hd__buf_1 _13190_ (.A(_06928_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_2 _13191_ (.A0(\core.cpuregs[20][16] ),
    .A1(_05377_),
    .S(_06922_),
    .X(_06929_));
 sky130_fd_sc_hd__buf_1 _13192_ (.A(_06929_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_2 _13193_ (.A0(\core.cpuregs[20][17] ),
    .A1(_05383_),
    .S(_06922_),
    .X(_06930_));
 sky130_fd_sc_hd__buf_1 _13194_ (.A(_06930_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_2 _13195_ (.A0(\core.cpuregs[20][18] ),
    .A1(_05388_),
    .S(_06922_),
    .X(_06931_));
 sky130_fd_sc_hd__buf_1 _13196_ (.A(_06931_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_2 _13197_ (.A0(\core.cpuregs[20][19] ),
    .A1(_05393_),
    .S(_06922_),
    .X(_06932_));
 sky130_fd_sc_hd__buf_1 _13198_ (.A(_06932_),
    .X(_00659_));
 sky130_fd_sc_hd__buf_1 _13199_ (.A(_06910_),
    .X(_06933_));
 sky130_fd_sc_hd__mux2_2 _13200_ (.A0(\core.cpuregs[20][20] ),
    .A1(_05399_),
    .S(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__buf_1 _13201_ (.A(_06934_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_2 _13202_ (.A0(\core.cpuregs[20][21] ),
    .A1(_05405_),
    .S(_06933_),
    .X(_06935_));
 sky130_fd_sc_hd__buf_1 _13203_ (.A(_06935_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_2 _13204_ (.A0(\core.cpuregs[20][22] ),
    .A1(_05410_),
    .S(_06933_),
    .X(_06936_));
 sky130_fd_sc_hd__buf_1 _13205_ (.A(_06936_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_2 _13206_ (.A0(\core.cpuregs[20][23] ),
    .A1(_05416_),
    .S(_06933_),
    .X(_06937_));
 sky130_fd_sc_hd__buf_1 _13207_ (.A(_06937_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_2 _13208_ (.A0(\core.cpuregs[20][24] ),
    .A1(_05421_),
    .S(_06933_),
    .X(_06938_));
 sky130_fd_sc_hd__buf_1 _13209_ (.A(_06938_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_2 _13210_ (.A0(\core.cpuregs[20][25] ),
    .A1(_05426_),
    .S(_06933_),
    .X(_06939_));
 sky130_fd_sc_hd__buf_1 _13211_ (.A(_06939_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_2 _13212_ (.A0(\core.cpuregs[20][26] ),
    .A1(_05432_),
    .S(_06933_),
    .X(_06940_));
 sky130_fd_sc_hd__buf_1 _13213_ (.A(_06940_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_2 _13214_ (.A0(\core.cpuregs[20][27] ),
    .A1(_05437_),
    .S(_06933_),
    .X(_06941_));
 sky130_fd_sc_hd__buf_1 _13215_ (.A(_06941_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_2 _13216_ (.A0(\core.cpuregs[20][28] ),
    .A1(_05442_),
    .S(_06933_),
    .X(_06942_));
 sky130_fd_sc_hd__buf_1 _13217_ (.A(_06942_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_2 _13218_ (.A0(\core.cpuregs[20][29] ),
    .A1(_05448_),
    .S(_06933_),
    .X(_06943_));
 sky130_fd_sc_hd__buf_1 _13219_ (.A(_06943_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_2 _13220_ (.A0(\core.cpuregs[20][30] ),
    .A1(_05453_),
    .S(_06910_),
    .X(_06944_));
 sky130_fd_sc_hd__buf_1 _13221_ (.A(_06944_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_2 _13222_ (.A0(\core.cpuregs[20][31] ),
    .A1(_05458_),
    .S(_06910_),
    .X(_06945_));
 sky130_fd_sc_hd__buf_1 _13223_ (.A(_06945_),
    .X(_00671_));
 sky130_fd_sc_hd__nor2_2 _13224_ (.A(_05657_),
    .B(_05837_),
    .Y(_06946_));
 sky130_fd_sc_hd__buf_1 _13225_ (.A(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__mux2_2 _13226_ (.A0(\core.cpuregs[25][0] ),
    .A1(_05284_),
    .S(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__buf_1 _13227_ (.A(_06948_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_2 _13228_ (.A0(\core.cpuregs[25][1] ),
    .A1(_05292_),
    .S(_06947_),
    .X(_06949_));
 sky130_fd_sc_hd__buf_1 _13229_ (.A(_06949_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_2 _13230_ (.A0(\core.cpuregs[25][2] ),
    .A1(_05297_),
    .S(_06947_),
    .X(_06950_));
 sky130_fd_sc_hd__buf_1 _13231_ (.A(_06950_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_2 _13232_ (.A0(\core.cpuregs[25][3] ),
    .A1(_05304_),
    .S(_06947_),
    .X(_06951_));
 sky130_fd_sc_hd__buf_1 _13233_ (.A(_06951_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_2 _13234_ (.A0(\core.cpuregs[25][4] ),
    .A1(_05310_),
    .S(_06947_),
    .X(_06952_));
 sky130_fd_sc_hd__buf_1 _13235_ (.A(_06952_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_2 _13236_ (.A0(\core.cpuregs[25][5] ),
    .A1(_05315_),
    .S(_06947_),
    .X(_06953_));
 sky130_fd_sc_hd__buf_1 _13237_ (.A(_06953_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_2 _13238_ (.A0(\core.cpuregs[25][6] ),
    .A1(_05320_),
    .S(_06947_),
    .X(_06954_));
 sky130_fd_sc_hd__buf_1 _13239_ (.A(_06954_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_2 _13240_ (.A0(\core.cpuregs[25][7] ),
    .A1(_05326_),
    .S(_06947_),
    .X(_06955_));
 sky130_fd_sc_hd__buf_1 _13241_ (.A(_06955_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_2 _13242_ (.A0(\core.cpuregs[25][8] ),
    .A1(_05332_),
    .S(_06947_),
    .X(_06956_));
 sky130_fd_sc_hd__buf_1 _13243_ (.A(_06956_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_2 _13244_ (.A0(\core.cpuregs[25][9] ),
    .A1(_05337_),
    .S(_06947_),
    .X(_06957_));
 sky130_fd_sc_hd__buf_1 _13245_ (.A(_06957_),
    .X(_00681_));
 sky130_fd_sc_hd__buf_1 _13246_ (.A(_06946_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_2 _13247_ (.A0(\core.cpuregs[25][10] ),
    .A1(_05343_),
    .S(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__buf_1 _13248_ (.A(_06959_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_2 _13249_ (.A0(\core.cpuregs[25][11] ),
    .A1(_05349_),
    .S(_06958_),
    .X(_06960_));
 sky130_fd_sc_hd__buf_1 _13250_ (.A(_06960_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_2 _13251_ (.A0(\core.cpuregs[25][12] ),
    .A1(_05355_),
    .S(_06958_),
    .X(_06961_));
 sky130_fd_sc_hd__buf_1 _13252_ (.A(_06961_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_2 _13253_ (.A0(\core.cpuregs[25][13] ),
    .A1(_05360_),
    .S(_06958_),
    .X(_06962_));
 sky130_fd_sc_hd__buf_1 _13254_ (.A(_06962_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_2 _13255_ (.A0(\core.cpuregs[25][14] ),
    .A1(_05367_),
    .S(_06958_),
    .X(_06963_));
 sky130_fd_sc_hd__buf_1 _13256_ (.A(_06963_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_2 _13257_ (.A0(\core.cpuregs[25][15] ),
    .A1(_05372_),
    .S(_06958_),
    .X(_06964_));
 sky130_fd_sc_hd__buf_1 _13258_ (.A(_06964_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_2 _13259_ (.A0(\core.cpuregs[25][16] ),
    .A1(_05377_),
    .S(_06958_),
    .X(_06965_));
 sky130_fd_sc_hd__buf_1 _13260_ (.A(_06965_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_2 _13261_ (.A0(\core.cpuregs[25][17] ),
    .A1(_05383_),
    .S(_06958_),
    .X(_06966_));
 sky130_fd_sc_hd__buf_1 _13262_ (.A(_06966_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_2 _13263_ (.A0(\core.cpuregs[25][18] ),
    .A1(_05388_),
    .S(_06958_),
    .X(_06967_));
 sky130_fd_sc_hd__buf_1 _13264_ (.A(_06967_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_2 _13265_ (.A0(\core.cpuregs[25][19] ),
    .A1(_05393_),
    .S(_06958_),
    .X(_06968_));
 sky130_fd_sc_hd__buf_1 _13266_ (.A(_06968_),
    .X(_00691_));
 sky130_fd_sc_hd__buf_1 _13267_ (.A(_06946_),
    .X(_06969_));
 sky130_fd_sc_hd__mux2_2 _13268_ (.A0(\core.cpuregs[25][20] ),
    .A1(_05399_),
    .S(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__buf_1 _13269_ (.A(_06970_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_2 _13270_ (.A0(\core.cpuregs[25][21] ),
    .A1(_05405_),
    .S(_06969_),
    .X(_06971_));
 sky130_fd_sc_hd__buf_1 _13271_ (.A(_06971_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_2 _13272_ (.A0(\core.cpuregs[25][22] ),
    .A1(_05410_),
    .S(_06969_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_1 _13273_ (.A(_06972_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_2 _13274_ (.A0(\core.cpuregs[25][23] ),
    .A1(_05416_),
    .S(_06969_),
    .X(_06973_));
 sky130_fd_sc_hd__buf_1 _13275_ (.A(_06973_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_2 _13276_ (.A0(\core.cpuregs[25][24] ),
    .A1(_05421_),
    .S(_06969_),
    .X(_06974_));
 sky130_fd_sc_hd__buf_1 _13277_ (.A(_06974_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_2 _13278_ (.A0(\core.cpuregs[25][25] ),
    .A1(_05426_),
    .S(_06969_),
    .X(_06975_));
 sky130_fd_sc_hd__buf_1 _13279_ (.A(_06975_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_2 _13280_ (.A0(\core.cpuregs[25][26] ),
    .A1(_05432_),
    .S(_06969_),
    .X(_06976_));
 sky130_fd_sc_hd__buf_1 _13281_ (.A(_06976_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_2 _13282_ (.A0(\core.cpuregs[25][27] ),
    .A1(_05437_),
    .S(_06969_),
    .X(_06977_));
 sky130_fd_sc_hd__buf_1 _13283_ (.A(_06977_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_2 _13284_ (.A0(\core.cpuregs[25][28] ),
    .A1(_05442_),
    .S(_06969_),
    .X(_06978_));
 sky130_fd_sc_hd__buf_1 _13285_ (.A(_06978_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_2 _13286_ (.A0(\core.cpuregs[25][29] ),
    .A1(_05448_),
    .S(_06969_),
    .X(_06979_));
 sky130_fd_sc_hd__buf_1 _13287_ (.A(_06979_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_2 _13288_ (.A0(\core.cpuregs[25][30] ),
    .A1(_05453_),
    .S(_06946_),
    .X(_06980_));
 sky130_fd_sc_hd__buf_1 _13289_ (.A(_06980_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_2 _13290_ (.A0(\core.cpuregs[25][31] ),
    .A1(_05458_),
    .S(_06946_),
    .X(_06981_));
 sky130_fd_sc_hd__buf_1 _13291_ (.A(_06981_),
    .X(_00703_));
 sky130_fd_sc_hd__or2_2 _13292_ (.A(_05620_),
    .B(_05837_),
    .X(_06982_));
 sky130_fd_sc_hd__buf_1 _13293_ (.A(_06982_),
    .X(_06983_));
 sky130_fd_sc_hd__mux2_2 _13294_ (.A0(_05460_),
    .A1(\core.cpuregs[1][0] ),
    .S(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__buf_1 _13295_ (.A(_06984_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_2 _13296_ (.A0(_05468_),
    .A1(\core.cpuregs[1][1] ),
    .S(_06983_),
    .X(_06985_));
 sky130_fd_sc_hd__buf_1 _13297_ (.A(_06985_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_2 _13298_ (.A0(_05470_),
    .A1(\core.cpuregs[1][2] ),
    .S(_06983_),
    .X(_06986_));
 sky130_fd_sc_hd__buf_1 _13299_ (.A(_06986_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_2 _13300_ (.A0(_05472_),
    .A1(\core.cpuregs[1][3] ),
    .S(_06983_),
    .X(_06987_));
 sky130_fd_sc_hd__buf_1 _13301_ (.A(_06987_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_2 _13302_ (.A0(_05474_),
    .A1(\core.cpuregs[1][4] ),
    .S(_06983_),
    .X(_06988_));
 sky130_fd_sc_hd__buf_1 _13303_ (.A(_06988_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_2 _13304_ (.A0(_05476_),
    .A1(\core.cpuregs[1][5] ),
    .S(_06983_),
    .X(_06989_));
 sky130_fd_sc_hd__buf_1 _13305_ (.A(_06989_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_2 _13306_ (.A0(_05478_),
    .A1(\core.cpuregs[1][6] ),
    .S(_06983_),
    .X(_06990_));
 sky130_fd_sc_hd__buf_1 _13307_ (.A(_06990_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_2 _13308_ (.A0(_05480_),
    .A1(\core.cpuregs[1][7] ),
    .S(_06983_),
    .X(_06991_));
 sky130_fd_sc_hd__buf_1 _13309_ (.A(_06991_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_2 _13310_ (.A0(_05482_),
    .A1(\core.cpuregs[1][8] ),
    .S(_06983_),
    .X(_06992_));
 sky130_fd_sc_hd__buf_1 _13311_ (.A(_06992_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_2 _13312_ (.A0(_05484_),
    .A1(\core.cpuregs[1][9] ),
    .S(_06983_),
    .X(_06993_));
 sky130_fd_sc_hd__buf_1 _13313_ (.A(_06993_),
    .X(_00713_));
 sky130_fd_sc_hd__buf_1 _13314_ (.A(_06982_),
    .X(_06994_));
 sky130_fd_sc_hd__mux2_2 _13315_ (.A0(_05486_),
    .A1(\core.cpuregs[1][10] ),
    .S(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__buf_1 _13316_ (.A(_06995_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_2 _13317_ (.A0(_05489_),
    .A1(\core.cpuregs[1][11] ),
    .S(_06994_),
    .X(_06996_));
 sky130_fd_sc_hd__buf_1 _13318_ (.A(_06996_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_2 _13319_ (.A0(_05491_),
    .A1(\core.cpuregs[1][12] ),
    .S(_06994_),
    .X(_06997_));
 sky130_fd_sc_hd__buf_1 _13320_ (.A(_06997_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_2 _13321_ (.A0(_05493_),
    .A1(\core.cpuregs[1][13] ),
    .S(_06994_),
    .X(_06998_));
 sky130_fd_sc_hd__buf_1 _13322_ (.A(_06998_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_2 _13323_ (.A0(_05495_),
    .A1(\core.cpuregs[1][14] ),
    .S(_06994_),
    .X(_06999_));
 sky130_fd_sc_hd__buf_1 _13324_ (.A(_06999_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_2 _13325_ (.A0(_05497_),
    .A1(\core.cpuregs[1][15] ),
    .S(_06994_),
    .X(_07000_));
 sky130_fd_sc_hd__buf_1 _13326_ (.A(_07000_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_2 _13327_ (.A0(_05499_),
    .A1(\core.cpuregs[1][16] ),
    .S(_06994_),
    .X(_07001_));
 sky130_fd_sc_hd__buf_1 _13328_ (.A(_07001_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_2 _13329_ (.A0(_05501_),
    .A1(\core.cpuregs[1][17] ),
    .S(_06994_),
    .X(_07002_));
 sky130_fd_sc_hd__buf_1 _13330_ (.A(_07002_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_2 _13331_ (.A0(_05503_),
    .A1(\core.cpuregs[1][18] ),
    .S(_06994_),
    .X(_07003_));
 sky130_fd_sc_hd__buf_1 _13332_ (.A(_07003_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_2 _13333_ (.A0(_05505_),
    .A1(\core.cpuregs[1][19] ),
    .S(_06994_),
    .X(_07004_));
 sky130_fd_sc_hd__buf_1 _13334_ (.A(_07004_),
    .X(_00723_));
 sky130_fd_sc_hd__buf_1 _13335_ (.A(_06982_),
    .X(_07005_));
 sky130_fd_sc_hd__mux2_2 _13336_ (.A0(_05507_),
    .A1(\core.cpuregs[1][20] ),
    .S(_07005_),
    .X(_07006_));
 sky130_fd_sc_hd__buf_1 _13337_ (.A(_07006_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_2 _13338_ (.A0(_05510_),
    .A1(\core.cpuregs[1][21] ),
    .S(_07005_),
    .X(_07007_));
 sky130_fd_sc_hd__buf_1 _13339_ (.A(_07007_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_2 _13340_ (.A0(_05512_),
    .A1(\core.cpuregs[1][22] ),
    .S(_07005_),
    .X(_07008_));
 sky130_fd_sc_hd__buf_1 _13341_ (.A(_07008_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_2 _13342_ (.A0(_05514_),
    .A1(\core.cpuregs[1][23] ),
    .S(_07005_),
    .X(_07009_));
 sky130_fd_sc_hd__buf_1 _13343_ (.A(_07009_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_2 _13344_ (.A0(_05516_),
    .A1(\core.cpuregs[1][24] ),
    .S(_07005_),
    .X(_07010_));
 sky130_fd_sc_hd__buf_1 _13345_ (.A(_07010_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_2 _13346_ (.A0(_05518_),
    .A1(\core.cpuregs[1][25] ),
    .S(_07005_),
    .X(_07011_));
 sky130_fd_sc_hd__buf_1 _13347_ (.A(_07011_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_2 _13348_ (.A0(_05520_),
    .A1(\core.cpuregs[1][26] ),
    .S(_07005_),
    .X(_07012_));
 sky130_fd_sc_hd__buf_1 _13349_ (.A(_07012_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_2 _13350_ (.A0(_05522_),
    .A1(\core.cpuregs[1][27] ),
    .S(_07005_),
    .X(_07013_));
 sky130_fd_sc_hd__buf_1 _13351_ (.A(_07013_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_2 _13352_ (.A0(_05524_),
    .A1(\core.cpuregs[1][28] ),
    .S(_07005_),
    .X(_07014_));
 sky130_fd_sc_hd__buf_1 _13353_ (.A(_07014_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_2 _13354_ (.A0(_05526_),
    .A1(\core.cpuregs[1][29] ),
    .S(_07005_),
    .X(_07015_));
 sky130_fd_sc_hd__buf_1 _13355_ (.A(_07015_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_2 _13356_ (.A0(_05528_),
    .A1(\core.cpuregs[1][30] ),
    .S(_06982_),
    .X(_07016_));
 sky130_fd_sc_hd__buf_1 _13357_ (.A(_07016_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_2 _13358_ (.A0(_05530_),
    .A1(\core.cpuregs[1][31] ),
    .S(_06982_),
    .X(_07017_));
 sky130_fd_sc_hd__buf_1 _13359_ (.A(_07017_),
    .X(_00735_));
 sky130_fd_sc_hd__buf_1 _13360_ (.A(_03176_),
    .X(_07018_));
 sky130_fd_sc_hd__mux2_2 _13361_ (.A0(\core.mem_rdata_q[7] ),
    .A1(mem_rdata[7]),
    .S(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__buf_1 _13362_ (.A(_07019_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_2 _13363_ (.A0(\core.decoded_rd[0] ),
    .A1(_01350_),
    .S(_03197_),
    .X(_07020_));
 sky130_fd_sc_hd__buf_1 _13364_ (.A(_07020_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_2 _13365_ (.A0(\core.mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(_07018_),
    .X(_07021_));
 sky130_fd_sc_hd__buf_1 _13366_ (.A(_07021_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_2 _13367_ (.A0(\core.decoded_rd[1] ),
    .A1(_01351_),
    .S(_03197_),
    .X(_07022_));
 sky130_fd_sc_hd__buf_1 _13368_ (.A(_07022_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_2 _13369_ (.A0(\core.mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(_07018_),
    .X(_07023_));
 sky130_fd_sc_hd__buf_1 _13370_ (.A(_07023_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_2 _13371_ (.A0(\core.decoded_rd[2] ),
    .A1(_01352_),
    .S(_03197_),
    .X(_07024_));
 sky130_fd_sc_hd__buf_1 _13372_ (.A(_07024_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_2 _13373_ (.A0(\core.mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(_07018_),
    .X(_07025_));
 sky130_fd_sc_hd__buf_1 _13374_ (.A(_07025_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_2 _13375_ (.A0(\core.decoded_rd[3] ),
    .A1(_01353_),
    .S(_03197_),
    .X(_07026_));
 sky130_fd_sc_hd__buf_1 _13376_ (.A(_07026_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_2 _13377_ (.A0(\core.mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(_07018_),
    .X(_07027_));
 sky130_fd_sc_hd__buf_1 _13378_ (.A(_07027_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_2 _13379_ (.A0(\core.decoded_rd[4] ),
    .A1(_01354_),
    .S(_03197_),
    .X(_07028_));
 sky130_fd_sc_hd__buf_1 _13380_ (.A(_07028_),
    .X(_00740_));
 sky130_fd_sc_hd__buf_1 _13381_ (.A(_05877_),
    .X(_07029_));
 sky130_fd_sc_hd__or3_2 _13382_ (.A(\core.instr_jalr ),
    .B(_02091_),
    .C(\core.is_alu_reg_imm ),
    .X(_07030_));
 sky130_fd_sc_hd__a221o_2 _13383_ (.A1(_02090_),
    .A2(\core.mem_rdata_q[7] ),
    .B1(\core.mem_rdata_q[20] ),
    .B2(_07030_),
    .C1(_05920_),
    .X(_07031_));
 sky130_fd_sc_hd__o21a_2 _13384_ (.A1(\core.decoded_imm[0] ),
    .A2(_07029_),
    .B1(_07031_),
    .X(_00741_));
 sky130_fd_sc_hd__buf_1 _13385_ (.A(_02448_),
    .X(_07032_));
 sky130_fd_sc_hd__mux2_2 _13386_ (.A0(\core.decoded_imm_j[1] ),
    .A1(_01364_),
    .S(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__buf_1 _13387_ (.A(_07033_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_2 _13388_ (.A0(\core.decoded_imm_j[2] ),
    .A1(_01365_),
    .S(_07032_),
    .X(_07034_));
 sky130_fd_sc_hd__buf_1 _13389_ (.A(_07034_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_2 _13390_ (.A0(\core.decoded_imm_j[3] ),
    .A1(_01366_),
    .S(_07032_),
    .X(_07035_));
 sky130_fd_sc_hd__buf_1 _13391_ (.A(_07035_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_2 _13392_ (.A0(\core.decoded_imm_j[4] ),
    .A1(_01367_),
    .S(_07032_),
    .X(_07036_));
 sky130_fd_sc_hd__buf_1 _13393_ (.A(_07036_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_2 _13394_ (.A0(\core.mem_rdata_q[25] ),
    .A1(mem_rdata[25]),
    .S(_07018_),
    .X(_07037_));
 sky130_fd_sc_hd__buf_1 _13395_ (.A(_07037_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_2 _13396_ (.A0(\core.decoded_imm_j[5] ),
    .A1(_01368_),
    .S(_03197_),
    .X(_07038_));
 sky130_fd_sc_hd__buf_1 _13397_ (.A(_07038_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_2 _13398_ (.A0(\core.mem_rdata_q[26] ),
    .A1(mem_rdata[26]),
    .S(_07018_),
    .X(_07039_));
 sky130_fd_sc_hd__buf_1 _13399_ (.A(_07039_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_2 _13400_ (.A0(\core.decoded_imm_j[6] ),
    .A1(_01369_),
    .S(_03197_),
    .X(_07040_));
 sky130_fd_sc_hd__buf_1 _13401_ (.A(_07040_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_2 _13402_ (.A0(\core.mem_rdata_q[27] ),
    .A1(mem_rdata[27]),
    .S(_07018_),
    .X(_07041_));
 sky130_fd_sc_hd__buf_1 _13403_ (.A(_07041_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_2 _13404_ (.A0(\core.decoded_imm_j[7] ),
    .A1(_01370_),
    .S(_03197_),
    .X(_07042_));
 sky130_fd_sc_hd__buf_1 _13405_ (.A(_07042_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_2 _13406_ (.A0(\core.mem_rdata_q[28] ),
    .A1(mem_rdata[28]),
    .S(_07018_),
    .X(_07043_));
 sky130_fd_sc_hd__buf_1 _13407_ (.A(_07043_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_2 _13408_ (.A0(\core.decoded_imm_j[8] ),
    .A1(_01371_),
    .S(_03197_),
    .X(_07044_));
 sky130_fd_sc_hd__buf_1 _13409_ (.A(_07044_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_2 _13410_ (.A0(\core.mem_rdata_q[29] ),
    .A1(mem_rdata[29]),
    .S(_07018_),
    .X(_07045_));
 sky130_fd_sc_hd__buf_1 _13411_ (.A(_07045_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_2 _13412_ (.A0(\core.decoded_imm_j[9] ),
    .A1(_01372_),
    .S(_07032_),
    .X(_07046_));
 sky130_fd_sc_hd__buf_1 _13413_ (.A(_07046_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_2 _13414_ (.A0(\core.mem_rdata_q[30] ),
    .A1(mem_rdata[30]),
    .S(_03177_),
    .X(_07047_));
 sky130_fd_sc_hd__buf_1 _13415_ (.A(_07047_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_2 _13416_ (.A0(\core.decoded_imm_j[10] ),
    .A1(_01373_),
    .S(_07032_),
    .X(_07048_));
 sky130_fd_sc_hd__buf_1 _13417_ (.A(_07048_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_2 _13418_ (.A0(\core.decoded_imm_j[11] ),
    .A1(_01363_),
    .S(_02448_),
    .X(_07049_));
 sky130_fd_sc_hd__buf_1 _13419_ (.A(_07049_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_2 _13420_ (.A0(\core.decoded_imm_j[12] ),
    .A1(_01355_),
    .S(_07032_),
    .X(_07050_));
 sky130_fd_sc_hd__buf_1 _13421_ (.A(_07050_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_2 _13422_ (.A0(\core.decoded_imm_j[13] ),
    .A1(_01356_),
    .S(_07032_),
    .X(_07051_));
 sky130_fd_sc_hd__buf_1 _13423_ (.A(_07051_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_2 _13424_ (.A0(\core.decoded_imm_j[14] ),
    .A1(_01357_),
    .S(_07032_),
    .X(_07052_));
 sky130_fd_sc_hd__buf_1 _13425_ (.A(_07052_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_2 _13426_ (.A0(\core.decoded_imm_j[15] ),
    .A1(_01358_),
    .S(_02448_),
    .X(_07053_));
 sky130_fd_sc_hd__buf_1 _13427_ (.A(_07053_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_2 _13428_ (.A0(\core.decoded_imm_j[16] ),
    .A1(_01359_),
    .S(_02448_),
    .X(_07054_));
 sky130_fd_sc_hd__buf_1 _13429_ (.A(_07054_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_2 _13430_ (.A0(\core.decoded_imm_j[17] ),
    .A1(_01360_),
    .S(_02448_),
    .X(_07055_));
 sky130_fd_sc_hd__buf_1 _13431_ (.A(_07055_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_2 _13432_ (.A0(\core.decoded_imm_j[18] ),
    .A1(_01361_),
    .S(_02448_),
    .X(_07056_));
 sky130_fd_sc_hd__buf_1 _13433_ (.A(_07056_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_2 _13434_ (.A0(\core.decoded_imm_j[19] ),
    .A1(_01362_),
    .S(_02448_),
    .X(_07057_));
 sky130_fd_sc_hd__buf_1 _13435_ (.A(_07057_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_2 _13436_ (.A0(\core.mem_rdata_q[31] ),
    .A1(mem_rdata[31]),
    .S(_03177_),
    .X(_07058_));
 sky130_fd_sc_hd__buf_1 _13437_ (.A(_07058_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_2 _13438_ (.A0(_04000_),
    .A1(_01374_),
    .S(_07032_),
    .X(_07059_));
 sky130_fd_sc_hd__buf_1 _13439_ (.A(_07059_),
    .X(_00761_));
 sky130_fd_sc_hd__nor2_2 _13440_ (.A(_01349_),
    .B(_01347_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_2 _13441_ (.A(_05814_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__a2bb2o_2 _13442_ (.A1_N(_01348_),
    .A2_N(_07061_),
    .B1(_02091_),
    .B2(_05803_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_2 _13443_ (.A(_05942_),
    .B(_05954_),
    .X(_07062_));
 sky130_fd_sc_hd__a22o_2 _13444_ (.A1(\core.is_slli_srli_srai ),
    .A2(_05921_),
    .B1(_05925_),
    .B2(_07062_),
    .X(_00763_));
 sky130_fd_sc_hd__a211o_2 _13445_ (.A1(\core.is_alu_reg_imm ),
    .A2(_05831_),
    .B1(_05943_),
    .C1(\core.instr_jalr ),
    .X(_07063_));
 sky130_fd_sc_hd__o21a_2 _13446_ (.A1(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ),
    .A2(_07029_),
    .B1(_07063_),
    .X(_00764_));
 sky130_fd_sc_hd__a32o_2 _13447_ (.A1(_01348_),
    .A2(_05814_),
    .A3(_07060_),
    .B1(_05803_),
    .B2(_02090_),
    .X(_00765_));
 sky130_fd_sc_hd__a22o_2 _13448_ (.A1(\core.is_sll_srl_sra ),
    .A2(_05921_),
    .B1(_05952_),
    .B2(_07062_),
    .X(_00766_));
 sky130_fd_sc_hd__a22o_2 _13449_ (.A1(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .A2(_05803_),
    .B1(_05814_),
    .B2(_05874_),
    .X(_07064_));
 sky130_fd_sc_hd__and2_2 _13450_ (.A(_05928_),
    .B(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__buf_1 _13451_ (.A(_07065_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_2 _13452_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .B(_02090_),
    .X(_07066_));
 sky130_fd_sc_hd__a221o_2 _13453_ (.A1(_03693_),
    .A2(_04000_),
    .B1(_07066_),
    .B2(\core.mem_rdata_q[31] ),
    .C1(_05830_),
    .X(_07067_));
 sky130_fd_sc_hd__buf_1 _13454_ (.A(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__buf_1 _13455_ (.A(_02020_),
    .X(_07069_));
 sky130_fd_sc_hd__o21a_2 _13456_ (.A1(_07069_),
    .A2(_07030_),
    .B1(\core.mem_rdata_q[31] ),
    .X(_07070_));
 sky130_fd_sc_hd__o22a_2 _13457_ (.A1(\core.decoded_imm[31] ),
    .A2(_07029_),
    .B1(_07068_),
    .B2(_07070_),
    .X(_00768_));
 sky130_fd_sc_hd__and2_2 _13458_ (.A(\core.mem_rdata_q[31] ),
    .B(_07030_),
    .X(_07071_));
 sky130_fd_sc_hd__buf_1 _13459_ (.A(_07071_),
    .X(_07072_));
 sky130_fd_sc_hd__a21o_2 _13460_ (.A1(\core.mem_rdata_q[30] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__o22a_2 _13461_ (.A1(\core.decoded_imm[30] ),
    .A2(_07029_),
    .B1(_07068_),
    .B2(_07073_),
    .X(_00769_));
 sky130_fd_sc_hd__buf_1 _13462_ (.A(_05877_),
    .X(_07074_));
 sky130_fd_sc_hd__a21o_2 _13463_ (.A1(\core.mem_rdata_q[29] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07075_));
 sky130_fd_sc_hd__o22a_2 _13464_ (.A1(\core.decoded_imm[29] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07075_),
    .X(_00770_));
 sky130_fd_sc_hd__a21o_2 _13465_ (.A1(\core.mem_rdata_q[28] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07076_));
 sky130_fd_sc_hd__o22a_2 _13466_ (.A1(\core.decoded_imm[28] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07076_),
    .X(_00771_));
 sky130_fd_sc_hd__a21o_2 _13467_ (.A1(\core.mem_rdata_q[27] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07077_));
 sky130_fd_sc_hd__o22a_2 _13468_ (.A1(\core.decoded_imm[27] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07077_),
    .X(_00772_));
 sky130_fd_sc_hd__a21o_2 _13469_ (.A1(\core.mem_rdata_q[26] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07078_));
 sky130_fd_sc_hd__o22a_2 _13470_ (.A1(\core.decoded_imm[26] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07078_),
    .X(_00773_));
 sky130_fd_sc_hd__a21o_2 _13471_ (.A1(\core.mem_rdata_q[25] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07079_));
 sky130_fd_sc_hd__o22a_2 _13472_ (.A1(\core.decoded_imm[25] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07079_),
    .X(_00774_));
 sky130_fd_sc_hd__a21o_2 _13473_ (.A1(\core.mem_rdata_q[24] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07080_));
 sky130_fd_sc_hd__o22a_2 _13474_ (.A1(\core.decoded_imm[24] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07080_),
    .X(_00775_));
 sky130_fd_sc_hd__a21o_2 _13475_ (.A1(\core.mem_rdata_q[23] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07081_));
 sky130_fd_sc_hd__o22a_2 _13476_ (.A1(\core.decoded_imm[23] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07081_),
    .X(_00776_));
 sky130_fd_sc_hd__a21o_2 _13477_ (.A1(\core.mem_rdata_q[22] ),
    .A2(_02021_),
    .B1(_07072_),
    .X(_07082_));
 sky130_fd_sc_hd__o22a_2 _13478_ (.A1(\core.decoded_imm[22] ),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07082_),
    .X(_00777_));
 sky130_fd_sc_hd__a21o_2 _13479_ (.A1(\core.mem_rdata_q[21] ),
    .A2(_07069_),
    .B1(_07072_),
    .X(_07083_));
 sky130_fd_sc_hd__o22a_2 _13480_ (.A1(\core.decoded_imm[21] ),
    .A2(_07074_),
    .B1(_07067_),
    .B2(_07083_),
    .X(_00778_));
 sky130_fd_sc_hd__a21o_2 _13481_ (.A1(\core.mem_rdata_q[20] ),
    .A2(_07069_),
    .B1(_07071_),
    .X(_07084_));
 sky130_fd_sc_hd__o22a_2 _13482_ (.A1(\core.decoded_imm[20] ),
    .A2(_07074_),
    .B1(_07067_),
    .B2(_07084_),
    .X(_00779_));
 sky130_fd_sc_hd__buf_1 _13483_ (.A(_05877_),
    .X(_07085_));
 sky130_fd_sc_hd__or3_2 _13484_ (.A(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .B(_02090_),
    .C(_07030_),
    .X(_07086_));
 sky130_fd_sc_hd__and2_2 _13485_ (.A(\core.mem_rdata_q[31] ),
    .B(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__buf_1 _13486_ (.A(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__buf_1 _13487_ (.A(_05830_),
    .X(_07089_));
 sky130_fd_sc_hd__a221o_2 _13488_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[19] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[19] ),
    .C1(_07089_),
    .X(_07090_));
 sky130_fd_sc_hd__o22a_2 _13489_ (.A1(\core.decoded_imm[19] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07090_),
    .X(_00780_));
 sky130_fd_sc_hd__a221o_2 _13490_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[18] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[18] ),
    .C1(_07089_),
    .X(_07091_));
 sky130_fd_sc_hd__o22a_2 _13491_ (.A1(\core.decoded_imm[18] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07091_),
    .X(_00781_));
 sky130_fd_sc_hd__buf_1 _13492_ (.A(_02018_),
    .X(_07092_));
 sky130_fd_sc_hd__a221o_2 _13493_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[17] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[17] ),
    .C1(_07089_),
    .X(_07093_));
 sky130_fd_sc_hd__o22a_2 _13494_ (.A1(\core.decoded_imm[17] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07093_),
    .X(_00782_));
 sky130_fd_sc_hd__a221o_2 _13495_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[16] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[16] ),
    .C1(_07089_),
    .X(_07094_));
 sky130_fd_sc_hd__o22a_2 _13496_ (.A1(\core.decoded_imm[16] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07094_),
    .X(_00783_));
 sky130_fd_sc_hd__a221o_2 _13497_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[15] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[15] ),
    .C1(_07089_),
    .X(_07095_));
 sky130_fd_sc_hd__o22a_2 _13498_ (.A1(\core.decoded_imm[15] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07095_),
    .X(_00784_));
 sky130_fd_sc_hd__a221o_2 _13499_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[14] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[14] ),
    .C1(_07089_),
    .X(_07096_));
 sky130_fd_sc_hd__o22a_2 _13500_ (.A1(\core.decoded_imm[14] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07096_),
    .X(_00785_));
 sky130_fd_sc_hd__a221o_2 _13501_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[13] ),
    .B1(_07069_),
    .B2(\core.mem_rdata_q[13] ),
    .C1(_07089_),
    .X(_07097_));
 sky130_fd_sc_hd__o22a_2 _13502_ (.A1(\core.decoded_imm[13] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07097_),
    .X(_00786_));
 sky130_fd_sc_hd__a221o_2 _13503_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[12] ),
    .B1(_02020_),
    .B2(\core.mem_rdata_q[12] ),
    .C1(_07089_),
    .X(_07098_));
 sky130_fd_sc_hd__o22a_2 _13504_ (.A1(\core.decoded_imm[12] ),
    .A2(_07085_),
    .B1(_07088_),
    .B2(_07098_),
    .X(_00787_));
 sky130_fd_sc_hd__o21a_2 _13505_ (.A1(_02090_),
    .A2(_07030_),
    .B1(\core.mem_rdata_q[31] ),
    .X(_07099_));
 sky130_fd_sc_hd__a221o_2 _13506_ (.A1(_02236_),
    .A2(\core.mem_rdata_q[7] ),
    .B1(\core.decoded_imm_j[11] ),
    .B2(_07092_),
    .C1(_07089_),
    .X(_07100_));
 sky130_fd_sc_hd__o22a_2 _13507_ (.A1(\core.decoded_imm[11] ),
    .A2(_07085_),
    .B1(_07099_),
    .B2(_07100_),
    .X(_00788_));
 sky130_fd_sc_hd__a221o_2 _13508_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[10] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[30] ),
    .C1(_05920_),
    .X(_07101_));
 sky130_fd_sc_hd__o21a_2 _13509_ (.A1(\core.decoded_imm[10] ),
    .A2(_07029_),
    .B1(_07101_),
    .X(_00789_));
 sky130_fd_sc_hd__a221o_2 _13510_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[9] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[29] ),
    .C1(_05920_),
    .X(_07102_));
 sky130_fd_sc_hd__o21a_2 _13511_ (.A1(\core.decoded_imm[9] ),
    .A2(_07029_),
    .B1(_07102_),
    .X(_00790_));
 sky130_fd_sc_hd__a221o_2 _13512_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[8] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[28] ),
    .C1(_05920_),
    .X(_07103_));
 sky130_fd_sc_hd__o21a_2 _13513_ (.A1(\core.decoded_imm[8] ),
    .A2(_07029_),
    .B1(_07103_),
    .X(_00791_));
 sky130_fd_sc_hd__a221o_2 _13514_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[7] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[27] ),
    .C1(_05920_),
    .X(_07104_));
 sky130_fd_sc_hd__o21a_2 _13515_ (.A1(\core.decoded_imm[7] ),
    .A2(_07029_),
    .B1(_07104_),
    .X(_00792_));
 sky130_fd_sc_hd__a221o_2 _13516_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[6] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[26] ),
    .C1(_05920_),
    .X(_07105_));
 sky130_fd_sc_hd__o21a_2 _13517_ (.A1(\core.decoded_imm[6] ),
    .A2(_07029_),
    .B1(_07105_),
    .X(_00793_));
 sky130_fd_sc_hd__a221o_2 _13518_ (.A1(_02019_),
    .A2(\core.decoded_imm_j[5] ),
    .B1(_07086_),
    .B2(\core.mem_rdata_q[25] ),
    .C1(_05920_),
    .X(_07106_));
 sky130_fd_sc_hd__o21a_2 _13519_ (.A1(\core.decoded_imm[5] ),
    .A2(_07029_),
    .B1(_07106_),
    .X(_00794_));
 sky130_fd_sc_hd__and2_2 _13520_ (.A(\core.mem_rdata_q[24] ),
    .B(_07030_),
    .X(_07107_));
 sky130_fd_sc_hd__a221o_2 _13521_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[4] ),
    .B1(_07066_),
    .B2(\core.mem_rdata_q[11] ),
    .C1(_05829_),
    .X(_07108_));
 sky130_fd_sc_hd__o22a_2 _13522_ (.A1(\core.decoded_imm[4] ),
    .A2(_07085_),
    .B1(_07107_),
    .B2(_07108_),
    .X(_00795_));
 sky130_fd_sc_hd__and2_2 _13523_ (.A(\core.mem_rdata_q[23] ),
    .B(_07030_),
    .X(_07109_));
 sky130_fd_sc_hd__a221o_2 _13524_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[3] ),
    .B1(_07066_),
    .B2(\core.mem_rdata_q[10] ),
    .C1(_05829_),
    .X(_07110_));
 sky130_fd_sc_hd__o22a_2 _13525_ (.A1(\core.decoded_imm[3] ),
    .A2(_05877_),
    .B1(_07109_),
    .B2(_07110_),
    .X(_00796_));
 sky130_fd_sc_hd__and2_2 _13526_ (.A(\core.mem_rdata_q[22] ),
    .B(_07030_),
    .X(_07111_));
 sky130_fd_sc_hd__a221o_2 _13527_ (.A1(_07092_),
    .A2(\core.decoded_imm_j[2] ),
    .B1(_07066_),
    .B2(\core.mem_rdata_q[9] ),
    .C1(_05829_),
    .X(_07112_));
 sky130_fd_sc_hd__o22a_2 _13528_ (.A1(\core.decoded_imm[2] ),
    .A2(_05877_),
    .B1(_07111_),
    .B2(_07112_),
    .X(_00797_));
 sky130_fd_sc_hd__a221o_2 _13529_ (.A1(\core.mem_rdata_q[21] ),
    .A2(_07030_),
    .B1(_07066_),
    .B2(\core.mem_rdata_q[8] ),
    .C1(_03660_),
    .X(_07113_));
 sky130_fd_sc_hd__mux2_2 _13530_ (.A0(\core.decoded_imm[1] ),
    .A1(_07113_),
    .S(_05877_),
    .X(_07114_));
 sky130_fd_sc_hd__buf_1 _13531_ (.A(_07114_),
    .X(_00798_));
 sky130_fd_sc_hd__or3b_2 _13532_ (.A(\core.latched_rd[3] ),
    .B(\core.latched_rd[2] ),
    .C_N(\core.latched_rd[4] ),
    .X(_07115_));
 sky130_fd_sc_hd__or2_2 _13533_ (.A(_05837_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__buf_1 _13534_ (.A(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__mux2_2 _13535_ (.A0(_05460_),
    .A1(\core.cpuregs[17][0] ),
    .S(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__buf_1 _13536_ (.A(_07118_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_2 _13537_ (.A0(_05468_),
    .A1(\core.cpuregs[17][1] ),
    .S(_07117_),
    .X(_07119_));
 sky130_fd_sc_hd__buf_1 _13538_ (.A(_07119_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_2 _13539_ (.A0(_05470_),
    .A1(\core.cpuregs[17][2] ),
    .S(_07117_),
    .X(_07120_));
 sky130_fd_sc_hd__buf_1 _13540_ (.A(_07120_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_2 _13541_ (.A0(_05472_),
    .A1(\core.cpuregs[17][3] ),
    .S(_07117_),
    .X(_07121_));
 sky130_fd_sc_hd__buf_1 _13542_ (.A(_07121_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_2 _13543_ (.A0(_05474_),
    .A1(\core.cpuregs[17][4] ),
    .S(_07117_),
    .X(_07122_));
 sky130_fd_sc_hd__buf_1 _13544_ (.A(_07122_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_2 _13545_ (.A0(_05476_),
    .A1(\core.cpuregs[17][5] ),
    .S(_07117_),
    .X(_07123_));
 sky130_fd_sc_hd__buf_1 _13546_ (.A(_07123_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_2 _13547_ (.A0(_05478_),
    .A1(\core.cpuregs[17][6] ),
    .S(_07117_),
    .X(_07124_));
 sky130_fd_sc_hd__buf_1 _13548_ (.A(_07124_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_2 _13549_ (.A0(_05480_),
    .A1(\core.cpuregs[17][7] ),
    .S(_07117_),
    .X(_07125_));
 sky130_fd_sc_hd__buf_1 _13550_ (.A(_07125_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_2 _13551_ (.A0(_05482_),
    .A1(\core.cpuregs[17][8] ),
    .S(_07117_),
    .X(_07126_));
 sky130_fd_sc_hd__buf_1 _13552_ (.A(_07126_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_2 _13553_ (.A0(_05484_),
    .A1(\core.cpuregs[17][9] ),
    .S(_07117_),
    .X(_07127_));
 sky130_fd_sc_hd__buf_1 _13554_ (.A(_07127_),
    .X(_00808_));
 sky130_fd_sc_hd__buf_1 _13555_ (.A(_07116_),
    .X(_07128_));
 sky130_fd_sc_hd__mux2_2 _13556_ (.A0(_05486_),
    .A1(\core.cpuregs[17][10] ),
    .S(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__buf_1 _13557_ (.A(_07129_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_2 _13558_ (.A0(_05489_),
    .A1(\core.cpuregs[17][11] ),
    .S(_07128_),
    .X(_07130_));
 sky130_fd_sc_hd__buf_1 _13559_ (.A(_07130_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_2 _13560_ (.A0(_05491_),
    .A1(\core.cpuregs[17][12] ),
    .S(_07128_),
    .X(_07131_));
 sky130_fd_sc_hd__buf_1 _13561_ (.A(_07131_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_2 _13562_ (.A0(_05493_),
    .A1(\core.cpuregs[17][13] ),
    .S(_07128_),
    .X(_07132_));
 sky130_fd_sc_hd__buf_1 _13563_ (.A(_07132_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_2 _13564_ (.A0(_05495_),
    .A1(\core.cpuregs[17][14] ),
    .S(_07128_),
    .X(_07133_));
 sky130_fd_sc_hd__buf_1 _13565_ (.A(_07133_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_2 _13566_ (.A0(_05497_),
    .A1(\core.cpuregs[17][15] ),
    .S(_07128_),
    .X(_07134_));
 sky130_fd_sc_hd__buf_1 _13567_ (.A(_07134_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_2 _13568_ (.A0(_05499_),
    .A1(\core.cpuregs[17][16] ),
    .S(_07128_),
    .X(_07135_));
 sky130_fd_sc_hd__buf_1 _13569_ (.A(_07135_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_2 _13570_ (.A0(_05501_),
    .A1(\core.cpuregs[17][17] ),
    .S(_07128_),
    .X(_07136_));
 sky130_fd_sc_hd__buf_1 _13571_ (.A(_07136_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_2 _13572_ (.A0(_05503_),
    .A1(\core.cpuregs[17][18] ),
    .S(_07128_),
    .X(_07137_));
 sky130_fd_sc_hd__buf_1 _13573_ (.A(_07137_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_2 _13574_ (.A0(_05505_),
    .A1(\core.cpuregs[17][19] ),
    .S(_07128_),
    .X(_07138_));
 sky130_fd_sc_hd__buf_1 _13575_ (.A(_07138_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_1 _13576_ (.A(_07116_),
    .X(_07139_));
 sky130_fd_sc_hd__mux2_2 _13577_ (.A0(_05507_),
    .A1(\core.cpuregs[17][20] ),
    .S(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__buf_1 _13578_ (.A(_07140_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_2 _13579_ (.A0(_05510_),
    .A1(\core.cpuregs[17][21] ),
    .S(_07139_),
    .X(_07141_));
 sky130_fd_sc_hd__buf_1 _13580_ (.A(_07141_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_2 _13581_ (.A0(_05512_),
    .A1(\core.cpuregs[17][22] ),
    .S(_07139_),
    .X(_07142_));
 sky130_fd_sc_hd__buf_1 _13582_ (.A(_07142_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_2 _13583_ (.A0(_05514_),
    .A1(\core.cpuregs[17][23] ),
    .S(_07139_),
    .X(_07143_));
 sky130_fd_sc_hd__buf_1 _13584_ (.A(_07143_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_2 _13585_ (.A0(_05516_),
    .A1(\core.cpuregs[17][24] ),
    .S(_07139_),
    .X(_07144_));
 sky130_fd_sc_hd__buf_1 _13586_ (.A(_07144_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_2 _13587_ (.A0(_05518_),
    .A1(\core.cpuregs[17][25] ),
    .S(_07139_),
    .X(_07145_));
 sky130_fd_sc_hd__buf_1 _13588_ (.A(_07145_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_2 _13589_ (.A0(_05520_),
    .A1(\core.cpuregs[17][26] ),
    .S(_07139_),
    .X(_07146_));
 sky130_fd_sc_hd__buf_1 _13590_ (.A(_07146_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_2 _13591_ (.A0(_05522_),
    .A1(\core.cpuregs[17][27] ),
    .S(_07139_),
    .X(_07147_));
 sky130_fd_sc_hd__buf_1 _13592_ (.A(_07147_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_2 _13593_ (.A0(_05524_),
    .A1(\core.cpuregs[17][28] ),
    .S(_07139_),
    .X(_07148_));
 sky130_fd_sc_hd__buf_1 _13594_ (.A(_07148_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_2 _13595_ (.A0(_05526_),
    .A1(\core.cpuregs[17][29] ),
    .S(_07139_),
    .X(_07149_));
 sky130_fd_sc_hd__buf_1 _13596_ (.A(_07149_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_2 _13597_ (.A0(_05528_),
    .A1(\core.cpuregs[17][30] ),
    .S(_07116_),
    .X(_07150_));
 sky130_fd_sc_hd__buf_1 _13598_ (.A(_07150_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_2 _13599_ (.A0(_05530_),
    .A1(\core.cpuregs[17][31] ),
    .S(_07116_),
    .X(_07151_));
 sky130_fd_sc_hd__buf_1 _13600_ (.A(_07151_),
    .X(_00830_));
 sky130_fd_sc_hd__or2_2 _13601_ (.A(_05766_),
    .B(_07115_),
    .X(_07152_));
 sky130_fd_sc_hd__buf_1 _13602_ (.A(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__mux2_2 _13603_ (.A0(_05460_),
    .A1(\core.cpuregs[16][0] ),
    .S(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__buf_1 _13604_ (.A(_07154_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_2 _13605_ (.A0(_05468_),
    .A1(\core.cpuregs[16][1] ),
    .S(_07153_),
    .X(_07155_));
 sky130_fd_sc_hd__buf_1 _13606_ (.A(_07155_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_2 _13607_ (.A0(_05470_),
    .A1(\core.cpuregs[16][2] ),
    .S(_07153_),
    .X(_07156_));
 sky130_fd_sc_hd__buf_1 _13608_ (.A(_07156_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_2 _13609_ (.A0(_05472_),
    .A1(\core.cpuregs[16][3] ),
    .S(_07153_),
    .X(_07157_));
 sky130_fd_sc_hd__buf_1 _13610_ (.A(_07157_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_2 _13611_ (.A0(_05474_),
    .A1(\core.cpuregs[16][4] ),
    .S(_07153_),
    .X(_07158_));
 sky130_fd_sc_hd__buf_1 _13612_ (.A(_07158_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_2 _13613_ (.A0(_05476_),
    .A1(\core.cpuregs[16][5] ),
    .S(_07153_),
    .X(_07159_));
 sky130_fd_sc_hd__buf_1 _13614_ (.A(_07159_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_2 _13615_ (.A0(_05478_),
    .A1(\core.cpuregs[16][6] ),
    .S(_07153_),
    .X(_07160_));
 sky130_fd_sc_hd__buf_1 _13616_ (.A(_07160_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_2 _13617_ (.A0(_05480_),
    .A1(\core.cpuregs[16][7] ),
    .S(_07153_),
    .X(_07161_));
 sky130_fd_sc_hd__buf_1 _13618_ (.A(_07161_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_2 _13619_ (.A0(_05482_),
    .A1(\core.cpuregs[16][8] ),
    .S(_07153_),
    .X(_07162_));
 sky130_fd_sc_hd__buf_1 _13620_ (.A(_07162_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_2 _13621_ (.A0(_05484_),
    .A1(\core.cpuregs[16][9] ),
    .S(_07153_),
    .X(_07163_));
 sky130_fd_sc_hd__buf_1 _13622_ (.A(_07163_),
    .X(_00840_));
 sky130_fd_sc_hd__buf_1 _13623_ (.A(_07152_),
    .X(_07164_));
 sky130_fd_sc_hd__mux2_2 _13624_ (.A0(_05486_),
    .A1(\core.cpuregs[16][10] ),
    .S(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__buf_1 _13625_ (.A(_07165_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_2 _13626_ (.A0(_05489_),
    .A1(\core.cpuregs[16][11] ),
    .S(_07164_),
    .X(_07166_));
 sky130_fd_sc_hd__buf_1 _13627_ (.A(_07166_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_2 _13628_ (.A0(_05491_),
    .A1(\core.cpuregs[16][12] ),
    .S(_07164_),
    .X(_07167_));
 sky130_fd_sc_hd__buf_1 _13629_ (.A(_07167_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_2 _13630_ (.A0(_05493_),
    .A1(\core.cpuregs[16][13] ),
    .S(_07164_),
    .X(_07168_));
 sky130_fd_sc_hd__buf_1 _13631_ (.A(_07168_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_2 _13632_ (.A0(_05495_),
    .A1(\core.cpuregs[16][14] ),
    .S(_07164_),
    .X(_07169_));
 sky130_fd_sc_hd__buf_1 _13633_ (.A(_07169_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_2 _13634_ (.A0(_05497_),
    .A1(\core.cpuregs[16][15] ),
    .S(_07164_),
    .X(_07170_));
 sky130_fd_sc_hd__buf_1 _13635_ (.A(_07170_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_2 _13636_ (.A0(_05499_),
    .A1(\core.cpuregs[16][16] ),
    .S(_07164_),
    .X(_07171_));
 sky130_fd_sc_hd__buf_1 _13637_ (.A(_07171_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_2 _13638_ (.A0(_05501_),
    .A1(\core.cpuregs[16][17] ),
    .S(_07164_),
    .X(_07172_));
 sky130_fd_sc_hd__buf_1 _13639_ (.A(_07172_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_2 _13640_ (.A0(_05503_),
    .A1(\core.cpuregs[16][18] ),
    .S(_07164_),
    .X(_07173_));
 sky130_fd_sc_hd__buf_1 _13641_ (.A(_07173_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_2 _13642_ (.A0(_05505_),
    .A1(\core.cpuregs[16][19] ),
    .S(_07164_),
    .X(_07174_));
 sky130_fd_sc_hd__buf_1 _13643_ (.A(_07174_),
    .X(_00850_));
 sky130_fd_sc_hd__buf_1 _13644_ (.A(_07152_),
    .X(_07175_));
 sky130_fd_sc_hd__mux2_2 _13645_ (.A0(_05507_),
    .A1(\core.cpuregs[16][20] ),
    .S(_07175_),
    .X(_07176_));
 sky130_fd_sc_hd__buf_1 _13646_ (.A(_07176_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_2 _13647_ (.A0(_05510_),
    .A1(\core.cpuregs[16][21] ),
    .S(_07175_),
    .X(_07177_));
 sky130_fd_sc_hd__buf_1 _13648_ (.A(_07177_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_2 _13649_ (.A0(_05512_),
    .A1(\core.cpuregs[16][22] ),
    .S(_07175_),
    .X(_07178_));
 sky130_fd_sc_hd__buf_1 _13650_ (.A(_07178_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_2 _13651_ (.A0(_05514_),
    .A1(\core.cpuregs[16][23] ),
    .S(_07175_),
    .X(_07179_));
 sky130_fd_sc_hd__buf_1 _13652_ (.A(_07179_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_2 _13653_ (.A0(_05516_),
    .A1(\core.cpuregs[16][24] ),
    .S(_07175_),
    .X(_07180_));
 sky130_fd_sc_hd__buf_1 _13654_ (.A(_07180_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_2 _13655_ (.A0(_05518_),
    .A1(\core.cpuregs[16][25] ),
    .S(_07175_),
    .X(_07181_));
 sky130_fd_sc_hd__buf_1 _13656_ (.A(_07181_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_2 _13657_ (.A0(_05520_),
    .A1(\core.cpuregs[16][26] ),
    .S(_07175_),
    .X(_07182_));
 sky130_fd_sc_hd__buf_1 _13658_ (.A(_07182_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_2 _13659_ (.A0(_05522_),
    .A1(\core.cpuregs[16][27] ),
    .S(_07175_),
    .X(_07183_));
 sky130_fd_sc_hd__buf_1 _13660_ (.A(_07183_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_2 _13661_ (.A0(_05524_),
    .A1(\core.cpuregs[16][28] ),
    .S(_07175_),
    .X(_07184_));
 sky130_fd_sc_hd__buf_1 _13662_ (.A(_07184_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_2 _13663_ (.A0(_05526_),
    .A1(\core.cpuregs[16][29] ),
    .S(_07175_),
    .X(_07185_));
 sky130_fd_sc_hd__buf_1 _13664_ (.A(_07185_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_2 _13665_ (.A0(_05528_),
    .A1(\core.cpuregs[16][30] ),
    .S(_07152_),
    .X(_07186_));
 sky130_fd_sc_hd__buf_1 _13666_ (.A(_07186_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_2 _13667_ (.A0(_05530_),
    .A1(\core.cpuregs[16][31] ),
    .S(_07152_),
    .X(_07187_));
 sky130_fd_sc_hd__buf_1 _13668_ (.A(_07187_),
    .X(_00862_));
 sky130_fd_sc_hd__buf_1 _13669_ (.A(_05283_),
    .X(_07188_));
 sky130_fd_sc_hd__nand3b_2 _13670_ (.A_N(\core.latched_rd[4] ),
    .B(\core.latched_rd[3] ),
    .C(\core.latched_rd[2] ),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_2 _13671_ (.A(_05286_),
    .B(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__buf_1 _13672_ (.A(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__mux2_2 _13673_ (.A0(\core.cpuregs[15][0] ),
    .A1(_07188_),
    .S(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__buf_1 _13674_ (.A(_07192_),
    .X(_00863_));
 sky130_fd_sc_hd__buf_1 _13675_ (.A(_05291_),
    .X(_07193_));
 sky130_fd_sc_hd__mux2_2 _13676_ (.A0(\core.cpuregs[15][1] ),
    .A1(_07193_),
    .S(_07191_),
    .X(_07194_));
 sky130_fd_sc_hd__buf_1 _13677_ (.A(_07194_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_1 _13678_ (.A(_05296_),
    .X(_07195_));
 sky130_fd_sc_hd__mux2_2 _13679_ (.A0(\core.cpuregs[15][2] ),
    .A1(_07195_),
    .S(_07191_),
    .X(_07196_));
 sky130_fd_sc_hd__buf_1 _13680_ (.A(_07196_),
    .X(_00865_));
 sky130_fd_sc_hd__buf_1 _13681_ (.A(_05303_),
    .X(_07197_));
 sky130_fd_sc_hd__mux2_2 _13682_ (.A0(\core.cpuregs[15][3] ),
    .A1(_07197_),
    .S(_07191_),
    .X(_07198_));
 sky130_fd_sc_hd__buf_1 _13683_ (.A(_07198_),
    .X(_00866_));
 sky130_fd_sc_hd__buf_1 _13684_ (.A(_05309_),
    .X(_07199_));
 sky130_fd_sc_hd__mux2_2 _13685_ (.A0(\core.cpuregs[15][4] ),
    .A1(_07199_),
    .S(_07191_),
    .X(_07200_));
 sky130_fd_sc_hd__buf_1 _13686_ (.A(_07200_),
    .X(_00867_));
 sky130_fd_sc_hd__buf_1 _13687_ (.A(_05314_),
    .X(_07201_));
 sky130_fd_sc_hd__mux2_2 _13688_ (.A0(\core.cpuregs[15][5] ),
    .A1(_07201_),
    .S(_07191_),
    .X(_07202_));
 sky130_fd_sc_hd__buf_1 _13689_ (.A(_07202_),
    .X(_00868_));
 sky130_fd_sc_hd__buf_1 _13690_ (.A(_05319_),
    .X(_07203_));
 sky130_fd_sc_hd__mux2_2 _13691_ (.A0(\core.cpuregs[15][6] ),
    .A1(_07203_),
    .S(_07191_),
    .X(_07204_));
 sky130_fd_sc_hd__buf_1 _13692_ (.A(_07204_),
    .X(_00869_));
 sky130_fd_sc_hd__buf_1 _13693_ (.A(_05325_),
    .X(_07205_));
 sky130_fd_sc_hd__mux2_2 _13694_ (.A0(\core.cpuregs[15][7] ),
    .A1(_07205_),
    .S(_07191_),
    .X(_07206_));
 sky130_fd_sc_hd__buf_1 _13695_ (.A(_07206_),
    .X(_00870_));
 sky130_fd_sc_hd__buf_1 _13696_ (.A(_05331_),
    .X(_07207_));
 sky130_fd_sc_hd__mux2_2 _13697_ (.A0(\core.cpuregs[15][8] ),
    .A1(_07207_),
    .S(_07191_),
    .X(_07208_));
 sky130_fd_sc_hd__buf_1 _13698_ (.A(_07208_),
    .X(_00871_));
 sky130_fd_sc_hd__buf_1 _13699_ (.A(_05336_),
    .X(_07209_));
 sky130_fd_sc_hd__mux2_2 _13700_ (.A0(\core.cpuregs[15][9] ),
    .A1(_07209_),
    .S(_07191_),
    .X(_07210_));
 sky130_fd_sc_hd__buf_1 _13701_ (.A(_07210_),
    .X(_00872_));
 sky130_fd_sc_hd__buf_1 _13702_ (.A(_05342_),
    .X(_07211_));
 sky130_fd_sc_hd__buf_1 _13703_ (.A(_07190_),
    .X(_07212_));
 sky130_fd_sc_hd__mux2_2 _13704_ (.A0(\core.cpuregs[15][10] ),
    .A1(_07211_),
    .S(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__buf_1 _13705_ (.A(_07213_),
    .X(_00873_));
 sky130_fd_sc_hd__buf_1 _13706_ (.A(_05348_),
    .X(_07214_));
 sky130_fd_sc_hd__mux2_2 _13707_ (.A0(\core.cpuregs[15][11] ),
    .A1(_07214_),
    .S(_07212_),
    .X(_07215_));
 sky130_fd_sc_hd__buf_1 _13708_ (.A(_07215_),
    .X(_00874_));
 sky130_fd_sc_hd__buf_1 _13709_ (.A(_05354_),
    .X(_07216_));
 sky130_fd_sc_hd__mux2_2 _13710_ (.A0(\core.cpuregs[15][12] ),
    .A1(_07216_),
    .S(_07212_),
    .X(_07217_));
 sky130_fd_sc_hd__buf_1 _13711_ (.A(_07217_),
    .X(_00875_));
 sky130_fd_sc_hd__buf_1 _13712_ (.A(_05359_),
    .X(_07218_));
 sky130_fd_sc_hd__mux2_2 _13713_ (.A0(\core.cpuregs[15][13] ),
    .A1(_07218_),
    .S(_07212_),
    .X(_07219_));
 sky130_fd_sc_hd__buf_1 _13714_ (.A(_07219_),
    .X(_00876_));
 sky130_fd_sc_hd__buf_1 _13715_ (.A(_05366_),
    .X(_07220_));
 sky130_fd_sc_hd__mux2_2 _13716_ (.A0(\core.cpuregs[15][14] ),
    .A1(_07220_),
    .S(_07212_),
    .X(_07221_));
 sky130_fd_sc_hd__buf_1 _13717_ (.A(_07221_),
    .X(_00877_));
 sky130_fd_sc_hd__buf_1 _13718_ (.A(_05371_),
    .X(_07222_));
 sky130_fd_sc_hd__mux2_2 _13719_ (.A0(\core.cpuregs[15][15] ),
    .A1(_07222_),
    .S(_07212_),
    .X(_07223_));
 sky130_fd_sc_hd__buf_1 _13720_ (.A(_07223_),
    .X(_00878_));
 sky130_fd_sc_hd__buf_1 _13721_ (.A(_05376_),
    .X(_07224_));
 sky130_fd_sc_hd__mux2_2 _13722_ (.A0(\core.cpuregs[15][16] ),
    .A1(_07224_),
    .S(_07212_),
    .X(_07225_));
 sky130_fd_sc_hd__buf_1 _13723_ (.A(_07225_),
    .X(_00879_));
 sky130_fd_sc_hd__buf_1 _13724_ (.A(_05382_),
    .X(_07226_));
 sky130_fd_sc_hd__mux2_2 _13725_ (.A0(\core.cpuregs[15][17] ),
    .A1(_07226_),
    .S(_07212_),
    .X(_07227_));
 sky130_fd_sc_hd__buf_1 _13726_ (.A(_07227_),
    .X(_00880_));
 sky130_fd_sc_hd__buf_1 _13727_ (.A(_05387_),
    .X(_07228_));
 sky130_fd_sc_hd__mux2_2 _13728_ (.A0(\core.cpuregs[15][18] ),
    .A1(_07228_),
    .S(_07212_),
    .X(_07229_));
 sky130_fd_sc_hd__buf_1 _13729_ (.A(_07229_),
    .X(_00881_));
 sky130_fd_sc_hd__buf_1 _13730_ (.A(_05392_),
    .X(_07230_));
 sky130_fd_sc_hd__mux2_2 _13731_ (.A0(\core.cpuregs[15][19] ),
    .A1(_07230_),
    .S(_07212_),
    .X(_07231_));
 sky130_fd_sc_hd__buf_1 _13732_ (.A(_07231_),
    .X(_00882_));
 sky130_fd_sc_hd__buf_1 _13733_ (.A(_05398_),
    .X(_07232_));
 sky130_fd_sc_hd__buf_1 _13734_ (.A(_07190_),
    .X(_07233_));
 sky130_fd_sc_hd__mux2_2 _13735_ (.A0(\core.cpuregs[15][20] ),
    .A1(_07232_),
    .S(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__buf_1 _13736_ (.A(_07234_),
    .X(_00883_));
 sky130_fd_sc_hd__buf_1 _13737_ (.A(_05404_),
    .X(_07235_));
 sky130_fd_sc_hd__mux2_2 _13738_ (.A0(\core.cpuregs[15][21] ),
    .A1(_07235_),
    .S(_07233_),
    .X(_07236_));
 sky130_fd_sc_hd__buf_1 _13739_ (.A(_07236_),
    .X(_00884_));
 sky130_fd_sc_hd__buf_1 _13740_ (.A(_05409_),
    .X(_07237_));
 sky130_fd_sc_hd__mux2_2 _13741_ (.A0(\core.cpuregs[15][22] ),
    .A1(_07237_),
    .S(_07233_),
    .X(_07238_));
 sky130_fd_sc_hd__buf_1 _13742_ (.A(_07238_),
    .X(_00885_));
 sky130_fd_sc_hd__buf_1 _13743_ (.A(_05415_),
    .X(_07239_));
 sky130_fd_sc_hd__mux2_2 _13744_ (.A0(\core.cpuregs[15][23] ),
    .A1(_07239_),
    .S(_07233_),
    .X(_07240_));
 sky130_fd_sc_hd__buf_1 _13745_ (.A(_07240_),
    .X(_00886_));
 sky130_fd_sc_hd__buf_1 _13746_ (.A(_05420_),
    .X(_07241_));
 sky130_fd_sc_hd__mux2_2 _13747_ (.A0(\core.cpuregs[15][24] ),
    .A1(_07241_),
    .S(_07233_),
    .X(_07242_));
 sky130_fd_sc_hd__buf_1 _13748_ (.A(_07242_),
    .X(_00887_));
 sky130_fd_sc_hd__buf_1 _13749_ (.A(_05425_),
    .X(_07243_));
 sky130_fd_sc_hd__mux2_2 _13750_ (.A0(\core.cpuregs[15][25] ),
    .A1(_07243_),
    .S(_07233_),
    .X(_07244_));
 sky130_fd_sc_hd__buf_1 _13751_ (.A(_07244_),
    .X(_00888_));
 sky130_fd_sc_hd__buf_1 _13752_ (.A(_05431_),
    .X(_07245_));
 sky130_fd_sc_hd__mux2_2 _13753_ (.A0(\core.cpuregs[15][26] ),
    .A1(_07245_),
    .S(_07233_),
    .X(_07246_));
 sky130_fd_sc_hd__buf_1 _13754_ (.A(_07246_),
    .X(_00889_));
 sky130_fd_sc_hd__buf_1 _13755_ (.A(_05436_),
    .X(_07247_));
 sky130_fd_sc_hd__mux2_2 _13756_ (.A0(\core.cpuregs[15][27] ),
    .A1(_07247_),
    .S(_07233_),
    .X(_07248_));
 sky130_fd_sc_hd__buf_1 _13757_ (.A(_07248_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_1 _13758_ (.A(_05441_),
    .X(_07249_));
 sky130_fd_sc_hd__mux2_2 _13759_ (.A0(\core.cpuregs[15][28] ),
    .A1(_07249_),
    .S(_07233_),
    .X(_07250_));
 sky130_fd_sc_hd__buf_1 _13760_ (.A(_07250_),
    .X(_00891_));
 sky130_fd_sc_hd__buf_1 _13761_ (.A(_05447_),
    .X(_07251_));
 sky130_fd_sc_hd__mux2_2 _13762_ (.A0(\core.cpuregs[15][29] ),
    .A1(_07251_),
    .S(_07233_),
    .X(_07252_));
 sky130_fd_sc_hd__buf_1 _13763_ (.A(_07252_),
    .X(_00892_));
 sky130_fd_sc_hd__buf_1 _13764_ (.A(_05452_),
    .X(_07253_));
 sky130_fd_sc_hd__mux2_2 _13765_ (.A0(\core.cpuregs[15][30] ),
    .A1(_07253_),
    .S(_07190_),
    .X(_07254_));
 sky130_fd_sc_hd__buf_1 _13766_ (.A(_07254_),
    .X(_00893_));
 sky130_fd_sc_hd__buf_1 _13767_ (.A(_05457_),
    .X(_07255_));
 sky130_fd_sc_hd__mux2_2 _13768_ (.A0(\core.cpuregs[15][31] ),
    .A1(_07255_),
    .S(_07190_),
    .X(_07256_));
 sky130_fd_sc_hd__buf_1 _13769_ (.A(_07256_),
    .X(_00894_));
 sky130_fd_sc_hd__or2_2 _13770_ (.A(_05464_),
    .B(_07189_),
    .X(_07257_));
 sky130_fd_sc_hd__buf_1 _13771_ (.A(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__mux2_2 _13772_ (.A0(_05460_),
    .A1(\core.cpuregs[14][0] ),
    .S(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__buf_1 _13773_ (.A(_07259_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_2 _13774_ (.A0(_05468_),
    .A1(\core.cpuregs[14][1] ),
    .S(_07258_),
    .X(_07260_));
 sky130_fd_sc_hd__buf_1 _13775_ (.A(_07260_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_2 _13776_ (.A0(_05470_),
    .A1(\core.cpuregs[14][2] ),
    .S(_07258_),
    .X(_07261_));
 sky130_fd_sc_hd__buf_1 _13777_ (.A(_07261_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_2 _13778_ (.A0(_05472_),
    .A1(\core.cpuregs[14][3] ),
    .S(_07258_),
    .X(_07262_));
 sky130_fd_sc_hd__buf_1 _13779_ (.A(_07262_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_2 _13780_ (.A0(_05474_),
    .A1(\core.cpuregs[14][4] ),
    .S(_07258_),
    .X(_07263_));
 sky130_fd_sc_hd__buf_1 _13781_ (.A(_07263_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_2 _13782_ (.A0(_05476_),
    .A1(\core.cpuregs[14][5] ),
    .S(_07258_),
    .X(_07264_));
 sky130_fd_sc_hd__buf_1 _13783_ (.A(_07264_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_2 _13784_ (.A0(_05478_),
    .A1(\core.cpuregs[14][6] ),
    .S(_07258_),
    .X(_07265_));
 sky130_fd_sc_hd__buf_1 _13785_ (.A(_07265_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_2 _13786_ (.A0(_05480_),
    .A1(\core.cpuregs[14][7] ),
    .S(_07258_),
    .X(_07266_));
 sky130_fd_sc_hd__buf_1 _13787_ (.A(_07266_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_2 _13788_ (.A0(_05482_),
    .A1(\core.cpuregs[14][8] ),
    .S(_07258_),
    .X(_07267_));
 sky130_fd_sc_hd__buf_1 _13789_ (.A(_07267_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_2 _13790_ (.A0(_05484_),
    .A1(\core.cpuregs[14][9] ),
    .S(_07258_),
    .X(_07268_));
 sky130_fd_sc_hd__buf_1 _13791_ (.A(_07268_),
    .X(_00904_));
 sky130_fd_sc_hd__buf_1 _13792_ (.A(_07257_),
    .X(_07269_));
 sky130_fd_sc_hd__mux2_2 _13793_ (.A0(_05486_),
    .A1(\core.cpuregs[14][10] ),
    .S(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__buf_1 _13794_ (.A(_07270_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_2 _13795_ (.A0(_05489_),
    .A1(\core.cpuregs[14][11] ),
    .S(_07269_),
    .X(_07271_));
 sky130_fd_sc_hd__buf_1 _13796_ (.A(_07271_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_2 _13797_ (.A0(_05491_),
    .A1(\core.cpuregs[14][12] ),
    .S(_07269_),
    .X(_07272_));
 sky130_fd_sc_hd__buf_1 _13798_ (.A(_07272_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_2 _13799_ (.A0(_05493_),
    .A1(\core.cpuregs[14][13] ),
    .S(_07269_),
    .X(_07273_));
 sky130_fd_sc_hd__buf_1 _13800_ (.A(_07273_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_2 _13801_ (.A0(_05495_),
    .A1(\core.cpuregs[14][14] ),
    .S(_07269_),
    .X(_07274_));
 sky130_fd_sc_hd__buf_1 _13802_ (.A(_07274_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_2 _13803_ (.A0(_05497_),
    .A1(\core.cpuregs[14][15] ),
    .S(_07269_),
    .X(_07275_));
 sky130_fd_sc_hd__buf_1 _13804_ (.A(_07275_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_2 _13805_ (.A0(_05499_),
    .A1(\core.cpuregs[14][16] ),
    .S(_07269_),
    .X(_07276_));
 sky130_fd_sc_hd__buf_1 _13806_ (.A(_07276_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_2 _13807_ (.A0(_05501_),
    .A1(\core.cpuregs[14][17] ),
    .S(_07269_),
    .X(_07277_));
 sky130_fd_sc_hd__buf_1 _13808_ (.A(_07277_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_2 _13809_ (.A0(_05503_),
    .A1(\core.cpuregs[14][18] ),
    .S(_07269_),
    .X(_07278_));
 sky130_fd_sc_hd__buf_1 _13810_ (.A(_07278_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_2 _13811_ (.A0(_05505_),
    .A1(\core.cpuregs[14][19] ),
    .S(_07269_),
    .X(_07279_));
 sky130_fd_sc_hd__buf_1 _13812_ (.A(_07279_),
    .X(_00914_));
 sky130_fd_sc_hd__buf_1 _13813_ (.A(_07257_),
    .X(_07280_));
 sky130_fd_sc_hd__mux2_2 _13814_ (.A0(_05507_),
    .A1(\core.cpuregs[14][20] ),
    .S(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__buf_1 _13815_ (.A(_07281_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_2 _13816_ (.A0(_05510_),
    .A1(\core.cpuregs[14][21] ),
    .S(_07280_),
    .X(_07282_));
 sky130_fd_sc_hd__buf_1 _13817_ (.A(_07282_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_2 _13818_ (.A0(_05512_),
    .A1(\core.cpuregs[14][22] ),
    .S(_07280_),
    .X(_07283_));
 sky130_fd_sc_hd__buf_1 _13819_ (.A(_07283_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_2 _13820_ (.A0(_05514_),
    .A1(\core.cpuregs[14][23] ),
    .S(_07280_),
    .X(_07284_));
 sky130_fd_sc_hd__buf_1 _13821_ (.A(_07284_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_2 _13822_ (.A0(_05516_),
    .A1(\core.cpuregs[14][24] ),
    .S(_07280_),
    .X(_07285_));
 sky130_fd_sc_hd__buf_1 _13823_ (.A(_07285_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_2 _13824_ (.A0(_05518_),
    .A1(\core.cpuregs[14][25] ),
    .S(_07280_),
    .X(_07286_));
 sky130_fd_sc_hd__buf_1 _13825_ (.A(_07286_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_2 _13826_ (.A0(_05520_),
    .A1(\core.cpuregs[14][26] ),
    .S(_07280_),
    .X(_07287_));
 sky130_fd_sc_hd__buf_1 _13827_ (.A(_07287_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_2 _13828_ (.A0(_05522_),
    .A1(\core.cpuregs[14][27] ),
    .S(_07280_),
    .X(_07288_));
 sky130_fd_sc_hd__buf_1 _13829_ (.A(_07288_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_2 _13830_ (.A0(_05524_),
    .A1(\core.cpuregs[14][28] ),
    .S(_07280_),
    .X(_07289_));
 sky130_fd_sc_hd__buf_1 _13831_ (.A(_07289_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_2 _13832_ (.A0(_05526_),
    .A1(\core.cpuregs[14][29] ),
    .S(_07280_),
    .X(_07290_));
 sky130_fd_sc_hd__buf_1 _13833_ (.A(_07290_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_2 _13834_ (.A0(_05528_),
    .A1(\core.cpuregs[14][30] ),
    .S(_07257_),
    .X(_07291_));
 sky130_fd_sc_hd__buf_1 _13835_ (.A(_07291_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_2 _13836_ (.A0(_05530_),
    .A1(\core.cpuregs[14][31] ),
    .S(_07257_),
    .X(_07292_));
 sky130_fd_sc_hd__buf_1 _13837_ (.A(_07292_),
    .X(_00926_));
 sky130_fd_sc_hd__nor2_2 _13838_ (.A(_05837_),
    .B(_07189_),
    .Y(_07293_));
 sky130_fd_sc_hd__buf_1 _13839_ (.A(_07293_),
    .X(_07294_));
 sky130_fd_sc_hd__mux2_2 _13840_ (.A0(\core.cpuregs[13][0] ),
    .A1(_07188_),
    .S(_07294_),
    .X(_07295_));
 sky130_fd_sc_hd__buf_1 _13841_ (.A(_07295_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_2 _13842_ (.A0(\core.cpuregs[13][1] ),
    .A1(_07193_),
    .S(_07294_),
    .X(_07296_));
 sky130_fd_sc_hd__buf_1 _13843_ (.A(_07296_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_2 _13844_ (.A0(\core.cpuregs[13][2] ),
    .A1(_07195_),
    .S(_07294_),
    .X(_07297_));
 sky130_fd_sc_hd__buf_1 _13845_ (.A(_07297_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_2 _13846_ (.A0(\core.cpuregs[13][3] ),
    .A1(_07197_),
    .S(_07294_),
    .X(_07298_));
 sky130_fd_sc_hd__buf_1 _13847_ (.A(_07298_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_2 _13848_ (.A0(\core.cpuregs[13][4] ),
    .A1(_07199_),
    .S(_07294_),
    .X(_07299_));
 sky130_fd_sc_hd__buf_1 _13849_ (.A(_07299_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_2 _13850_ (.A0(\core.cpuregs[13][5] ),
    .A1(_07201_),
    .S(_07294_),
    .X(_07300_));
 sky130_fd_sc_hd__buf_1 _13851_ (.A(_07300_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_2 _13852_ (.A0(\core.cpuregs[13][6] ),
    .A1(_07203_),
    .S(_07294_),
    .X(_07301_));
 sky130_fd_sc_hd__buf_1 _13853_ (.A(_07301_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_2 _13854_ (.A0(\core.cpuregs[13][7] ),
    .A1(_07205_),
    .S(_07294_),
    .X(_07302_));
 sky130_fd_sc_hd__buf_1 _13855_ (.A(_07302_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_2 _13856_ (.A0(\core.cpuregs[13][8] ),
    .A1(_07207_),
    .S(_07294_),
    .X(_07303_));
 sky130_fd_sc_hd__buf_1 _13857_ (.A(_07303_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_2 _13858_ (.A0(\core.cpuregs[13][9] ),
    .A1(_07209_),
    .S(_07294_),
    .X(_07304_));
 sky130_fd_sc_hd__buf_1 _13859_ (.A(_07304_),
    .X(_00936_));
 sky130_fd_sc_hd__buf_1 _13860_ (.A(_07293_),
    .X(_07305_));
 sky130_fd_sc_hd__mux2_2 _13861_ (.A0(\core.cpuregs[13][10] ),
    .A1(_07211_),
    .S(_07305_),
    .X(_07306_));
 sky130_fd_sc_hd__buf_1 _13862_ (.A(_07306_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_2 _13863_ (.A0(\core.cpuregs[13][11] ),
    .A1(_07214_),
    .S(_07305_),
    .X(_07307_));
 sky130_fd_sc_hd__buf_1 _13864_ (.A(_07307_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_2 _13865_ (.A0(\core.cpuregs[13][12] ),
    .A1(_07216_),
    .S(_07305_),
    .X(_07308_));
 sky130_fd_sc_hd__buf_1 _13866_ (.A(_07308_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_2 _13867_ (.A0(\core.cpuregs[13][13] ),
    .A1(_07218_),
    .S(_07305_),
    .X(_07309_));
 sky130_fd_sc_hd__buf_1 _13868_ (.A(_07309_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_2 _13869_ (.A0(\core.cpuregs[13][14] ),
    .A1(_07220_),
    .S(_07305_),
    .X(_07310_));
 sky130_fd_sc_hd__buf_1 _13870_ (.A(_07310_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_2 _13871_ (.A0(\core.cpuregs[13][15] ),
    .A1(_07222_),
    .S(_07305_),
    .X(_07311_));
 sky130_fd_sc_hd__buf_1 _13872_ (.A(_07311_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_2 _13873_ (.A0(\core.cpuregs[13][16] ),
    .A1(_07224_),
    .S(_07305_),
    .X(_07312_));
 sky130_fd_sc_hd__buf_1 _13874_ (.A(_07312_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_2 _13875_ (.A0(\core.cpuregs[13][17] ),
    .A1(_07226_),
    .S(_07305_),
    .X(_07313_));
 sky130_fd_sc_hd__buf_1 _13876_ (.A(_07313_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_2 _13877_ (.A0(\core.cpuregs[13][18] ),
    .A1(_07228_),
    .S(_07305_),
    .X(_07314_));
 sky130_fd_sc_hd__buf_1 _13878_ (.A(_07314_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_2 _13879_ (.A0(\core.cpuregs[13][19] ),
    .A1(_07230_),
    .S(_07305_),
    .X(_07315_));
 sky130_fd_sc_hd__buf_1 _13880_ (.A(_07315_),
    .X(_00946_));
 sky130_fd_sc_hd__buf_1 _13881_ (.A(_07293_),
    .X(_07316_));
 sky130_fd_sc_hd__mux2_2 _13882_ (.A0(\core.cpuregs[13][20] ),
    .A1(_07232_),
    .S(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__buf_1 _13883_ (.A(_07317_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_2 _13884_ (.A0(\core.cpuregs[13][21] ),
    .A1(_07235_),
    .S(_07316_),
    .X(_07318_));
 sky130_fd_sc_hd__buf_1 _13885_ (.A(_07318_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_2 _13886_ (.A0(\core.cpuregs[13][22] ),
    .A1(_07237_),
    .S(_07316_),
    .X(_07319_));
 sky130_fd_sc_hd__buf_1 _13887_ (.A(_07319_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_2 _13888_ (.A0(\core.cpuregs[13][23] ),
    .A1(_07239_),
    .S(_07316_),
    .X(_07320_));
 sky130_fd_sc_hd__buf_1 _13889_ (.A(_07320_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_2 _13890_ (.A0(\core.cpuregs[13][24] ),
    .A1(_07241_),
    .S(_07316_),
    .X(_07321_));
 sky130_fd_sc_hd__buf_1 _13891_ (.A(_07321_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_2 _13892_ (.A0(\core.cpuregs[13][25] ),
    .A1(_07243_),
    .S(_07316_),
    .X(_07322_));
 sky130_fd_sc_hd__buf_1 _13893_ (.A(_07322_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_2 _13894_ (.A0(\core.cpuregs[13][26] ),
    .A1(_07245_),
    .S(_07316_),
    .X(_07323_));
 sky130_fd_sc_hd__buf_1 _13895_ (.A(_07323_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_2 _13896_ (.A0(\core.cpuregs[13][27] ),
    .A1(_07247_),
    .S(_07316_),
    .X(_07324_));
 sky130_fd_sc_hd__buf_1 _13897_ (.A(_07324_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_2 _13898_ (.A0(\core.cpuregs[13][28] ),
    .A1(_07249_),
    .S(_07316_),
    .X(_07325_));
 sky130_fd_sc_hd__buf_1 _13899_ (.A(_07325_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_2 _13900_ (.A0(\core.cpuregs[13][29] ),
    .A1(_07251_),
    .S(_07316_),
    .X(_07326_));
 sky130_fd_sc_hd__buf_1 _13901_ (.A(_07326_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_2 _13902_ (.A0(\core.cpuregs[13][30] ),
    .A1(_07253_),
    .S(_07293_),
    .X(_07327_));
 sky130_fd_sc_hd__buf_1 _13903_ (.A(_07327_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_2 _13904_ (.A0(\core.cpuregs[13][31] ),
    .A1(_07255_),
    .S(_07293_),
    .X(_07328_));
 sky130_fd_sc_hd__buf_1 _13905_ (.A(_07328_),
    .X(_00958_));
 sky130_fd_sc_hd__nor2_2 _13906_ (.A(_05766_),
    .B(_07189_),
    .Y(_07329_));
 sky130_fd_sc_hd__buf_1 _13907_ (.A(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__mux2_2 _13908_ (.A0(\core.cpuregs[12][0] ),
    .A1(_07188_),
    .S(_07330_),
    .X(_07331_));
 sky130_fd_sc_hd__buf_1 _13909_ (.A(_07331_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_2 _13910_ (.A0(\core.cpuregs[12][1] ),
    .A1(_07193_),
    .S(_07330_),
    .X(_07332_));
 sky130_fd_sc_hd__buf_1 _13911_ (.A(_07332_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_2 _13912_ (.A0(\core.cpuregs[12][2] ),
    .A1(_07195_),
    .S(_07330_),
    .X(_07333_));
 sky130_fd_sc_hd__buf_1 _13913_ (.A(_07333_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_2 _13914_ (.A0(\core.cpuregs[12][3] ),
    .A1(_07197_),
    .S(_07330_),
    .X(_07334_));
 sky130_fd_sc_hd__buf_1 _13915_ (.A(_07334_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_2 _13916_ (.A0(\core.cpuregs[12][4] ),
    .A1(_07199_),
    .S(_07330_),
    .X(_07335_));
 sky130_fd_sc_hd__buf_1 _13917_ (.A(_07335_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_2 _13918_ (.A0(\core.cpuregs[12][5] ),
    .A1(_07201_),
    .S(_07330_),
    .X(_07336_));
 sky130_fd_sc_hd__buf_1 _13919_ (.A(_07336_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_2 _13920_ (.A0(\core.cpuregs[12][6] ),
    .A1(_07203_),
    .S(_07330_),
    .X(_07337_));
 sky130_fd_sc_hd__buf_1 _13921_ (.A(_07337_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_2 _13922_ (.A0(\core.cpuregs[12][7] ),
    .A1(_07205_),
    .S(_07330_),
    .X(_07338_));
 sky130_fd_sc_hd__buf_1 _13923_ (.A(_07338_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_2 _13924_ (.A0(\core.cpuregs[12][8] ),
    .A1(_07207_),
    .S(_07330_),
    .X(_07339_));
 sky130_fd_sc_hd__buf_1 _13925_ (.A(_07339_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_2 _13926_ (.A0(\core.cpuregs[12][9] ),
    .A1(_07209_),
    .S(_07330_),
    .X(_07340_));
 sky130_fd_sc_hd__buf_1 _13927_ (.A(_07340_),
    .X(_00968_));
 sky130_fd_sc_hd__buf_1 _13928_ (.A(_07329_),
    .X(_07341_));
 sky130_fd_sc_hd__mux2_2 _13929_ (.A0(\core.cpuregs[12][10] ),
    .A1(_07211_),
    .S(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__buf_1 _13930_ (.A(_07342_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_2 _13931_ (.A0(\core.cpuregs[12][11] ),
    .A1(_07214_),
    .S(_07341_),
    .X(_07343_));
 sky130_fd_sc_hd__buf_1 _13932_ (.A(_07343_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_2 _13933_ (.A0(\core.cpuregs[12][12] ),
    .A1(_07216_),
    .S(_07341_),
    .X(_07344_));
 sky130_fd_sc_hd__buf_1 _13934_ (.A(_07344_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_2 _13935_ (.A0(\core.cpuregs[12][13] ),
    .A1(_07218_),
    .S(_07341_),
    .X(_07345_));
 sky130_fd_sc_hd__buf_1 _13936_ (.A(_07345_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_2 _13937_ (.A0(\core.cpuregs[12][14] ),
    .A1(_07220_),
    .S(_07341_),
    .X(_07346_));
 sky130_fd_sc_hd__buf_1 _13938_ (.A(_07346_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_2 _13939_ (.A0(\core.cpuregs[12][15] ),
    .A1(_07222_),
    .S(_07341_),
    .X(_07347_));
 sky130_fd_sc_hd__buf_1 _13940_ (.A(_07347_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_2 _13941_ (.A0(\core.cpuregs[12][16] ),
    .A1(_07224_),
    .S(_07341_),
    .X(_07348_));
 sky130_fd_sc_hd__buf_1 _13942_ (.A(_07348_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_2 _13943_ (.A0(\core.cpuregs[12][17] ),
    .A1(_07226_),
    .S(_07341_),
    .X(_07349_));
 sky130_fd_sc_hd__buf_1 _13944_ (.A(_07349_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_2 _13945_ (.A0(\core.cpuregs[12][18] ),
    .A1(_07228_),
    .S(_07341_),
    .X(_07350_));
 sky130_fd_sc_hd__buf_1 _13946_ (.A(_07350_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_2 _13947_ (.A0(\core.cpuregs[12][19] ),
    .A1(_07230_),
    .S(_07341_),
    .X(_07351_));
 sky130_fd_sc_hd__buf_1 _13948_ (.A(_07351_),
    .X(_00978_));
 sky130_fd_sc_hd__buf_1 _13949_ (.A(_07329_),
    .X(_07352_));
 sky130_fd_sc_hd__mux2_2 _13950_ (.A0(\core.cpuregs[12][20] ),
    .A1(_07232_),
    .S(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__buf_1 _13951_ (.A(_07353_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_2 _13952_ (.A0(\core.cpuregs[12][21] ),
    .A1(_07235_),
    .S(_07352_),
    .X(_07354_));
 sky130_fd_sc_hd__buf_1 _13953_ (.A(_07354_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_2 _13954_ (.A0(\core.cpuregs[12][22] ),
    .A1(_07237_),
    .S(_07352_),
    .X(_07355_));
 sky130_fd_sc_hd__buf_1 _13955_ (.A(_07355_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_2 _13956_ (.A0(\core.cpuregs[12][23] ),
    .A1(_07239_),
    .S(_07352_),
    .X(_07356_));
 sky130_fd_sc_hd__buf_1 _13957_ (.A(_07356_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_2 _13958_ (.A0(\core.cpuregs[12][24] ),
    .A1(_07241_),
    .S(_07352_),
    .X(_07357_));
 sky130_fd_sc_hd__buf_1 _13959_ (.A(_07357_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_2 _13960_ (.A0(\core.cpuregs[12][25] ),
    .A1(_07243_),
    .S(_07352_),
    .X(_07358_));
 sky130_fd_sc_hd__buf_1 _13961_ (.A(_07358_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_2 _13962_ (.A0(\core.cpuregs[12][26] ),
    .A1(_07245_),
    .S(_07352_),
    .X(_07359_));
 sky130_fd_sc_hd__buf_1 _13963_ (.A(_07359_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_2 _13964_ (.A0(\core.cpuregs[12][27] ),
    .A1(_07247_),
    .S(_07352_),
    .X(_07360_));
 sky130_fd_sc_hd__buf_1 _13965_ (.A(_07360_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_2 _13966_ (.A0(\core.cpuregs[12][28] ),
    .A1(_07249_),
    .S(_07352_),
    .X(_07361_));
 sky130_fd_sc_hd__buf_1 _13967_ (.A(_07361_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_2 _13968_ (.A0(\core.cpuregs[12][29] ),
    .A1(_07251_),
    .S(_07352_),
    .X(_07362_));
 sky130_fd_sc_hd__buf_1 _13969_ (.A(_07362_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_2 _13970_ (.A0(\core.cpuregs[12][30] ),
    .A1(_07253_),
    .S(_07329_),
    .X(_07363_));
 sky130_fd_sc_hd__buf_1 _13971_ (.A(_07363_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_2 _13972_ (.A0(\core.cpuregs[12][31] ),
    .A1(_07255_),
    .S(_07329_),
    .X(_07364_));
 sky130_fd_sc_hd__buf_1 _13973_ (.A(_07364_),
    .X(_00990_));
 sky130_fd_sc_hd__or3b_2 _13974_ (.A(\core.latched_rd[4] ),
    .B(\core.latched_rd[2] ),
    .C_N(\core.latched_rd[3] ),
    .X(_07365_));
 sky130_fd_sc_hd__nor2_2 _13975_ (.A(_05286_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__buf_1 _13976_ (.A(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__mux2_2 _13977_ (.A0(\core.cpuregs[11][0] ),
    .A1(_07188_),
    .S(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__buf_1 _13978_ (.A(_07368_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_2 _13979_ (.A0(\core.cpuregs[11][1] ),
    .A1(_07193_),
    .S(_07367_),
    .X(_07369_));
 sky130_fd_sc_hd__buf_1 _13980_ (.A(_07369_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_2 _13981_ (.A0(\core.cpuregs[11][2] ),
    .A1(_07195_),
    .S(_07367_),
    .X(_07370_));
 sky130_fd_sc_hd__buf_1 _13982_ (.A(_07370_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_2 _13983_ (.A0(\core.cpuregs[11][3] ),
    .A1(_07197_),
    .S(_07367_),
    .X(_07371_));
 sky130_fd_sc_hd__buf_1 _13984_ (.A(_07371_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_2 _13985_ (.A0(\core.cpuregs[11][4] ),
    .A1(_07199_),
    .S(_07367_),
    .X(_07372_));
 sky130_fd_sc_hd__buf_1 _13986_ (.A(_07372_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_2 _13987_ (.A0(\core.cpuregs[11][5] ),
    .A1(_07201_),
    .S(_07367_),
    .X(_07373_));
 sky130_fd_sc_hd__buf_1 _13988_ (.A(_07373_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_2 _13989_ (.A0(\core.cpuregs[11][6] ),
    .A1(_07203_),
    .S(_07367_),
    .X(_07374_));
 sky130_fd_sc_hd__buf_1 _13990_ (.A(_07374_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_2 _13991_ (.A0(\core.cpuregs[11][7] ),
    .A1(_07205_),
    .S(_07367_),
    .X(_07375_));
 sky130_fd_sc_hd__buf_1 _13992_ (.A(_07375_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_2 _13993_ (.A0(\core.cpuregs[11][8] ),
    .A1(_07207_),
    .S(_07367_),
    .X(_07376_));
 sky130_fd_sc_hd__buf_1 _13994_ (.A(_07376_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_2 _13995_ (.A0(\core.cpuregs[11][9] ),
    .A1(_07209_),
    .S(_07367_),
    .X(_07377_));
 sky130_fd_sc_hd__buf_1 _13996_ (.A(_07377_),
    .X(_01000_));
 sky130_fd_sc_hd__buf_1 _13997_ (.A(_07366_),
    .X(_07378_));
 sky130_fd_sc_hd__mux2_2 _13998_ (.A0(\core.cpuregs[11][10] ),
    .A1(_07211_),
    .S(_07378_),
    .X(_07379_));
 sky130_fd_sc_hd__buf_1 _13999_ (.A(_07379_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_2 _14000_ (.A0(\core.cpuregs[11][11] ),
    .A1(_07214_),
    .S(_07378_),
    .X(_07380_));
 sky130_fd_sc_hd__buf_1 _14001_ (.A(_07380_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_2 _14002_ (.A0(\core.cpuregs[11][12] ),
    .A1(_07216_),
    .S(_07378_),
    .X(_07381_));
 sky130_fd_sc_hd__buf_1 _14003_ (.A(_07381_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_2 _14004_ (.A0(\core.cpuregs[11][13] ),
    .A1(_07218_),
    .S(_07378_),
    .X(_07382_));
 sky130_fd_sc_hd__buf_1 _14005_ (.A(_07382_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_2 _14006_ (.A0(\core.cpuregs[11][14] ),
    .A1(_07220_),
    .S(_07378_),
    .X(_07383_));
 sky130_fd_sc_hd__buf_1 _14007_ (.A(_07383_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_2 _14008_ (.A0(\core.cpuregs[11][15] ),
    .A1(_07222_),
    .S(_07378_),
    .X(_07384_));
 sky130_fd_sc_hd__buf_1 _14009_ (.A(_07384_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_2 _14010_ (.A0(\core.cpuregs[11][16] ),
    .A1(_07224_),
    .S(_07378_),
    .X(_07385_));
 sky130_fd_sc_hd__buf_1 _14011_ (.A(_07385_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_2 _14012_ (.A0(\core.cpuregs[11][17] ),
    .A1(_07226_),
    .S(_07378_),
    .X(_07386_));
 sky130_fd_sc_hd__buf_1 _14013_ (.A(_07386_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_2 _14014_ (.A0(\core.cpuregs[11][18] ),
    .A1(_07228_),
    .S(_07378_),
    .X(_07387_));
 sky130_fd_sc_hd__buf_1 _14015_ (.A(_07387_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_2 _14016_ (.A0(\core.cpuregs[11][19] ),
    .A1(_07230_),
    .S(_07378_),
    .X(_07388_));
 sky130_fd_sc_hd__buf_1 _14017_ (.A(_07388_),
    .X(_01010_));
 sky130_fd_sc_hd__buf_1 _14018_ (.A(_07366_),
    .X(_07389_));
 sky130_fd_sc_hd__mux2_2 _14019_ (.A0(\core.cpuregs[11][20] ),
    .A1(_07232_),
    .S(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__buf_1 _14020_ (.A(_07390_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_2 _14021_ (.A0(\core.cpuregs[11][21] ),
    .A1(_07235_),
    .S(_07389_),
    .X(_07391_));
 sky130_fd_sc_hd__buf_1 _14022_ (.A(_07391_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_2 _14023_ (.A0(\core.cpuregs[11][22] ),
    .A1(_07237_),
    .S(_07389_),
    .X(_07392_));
 sky130_fd_sc_hd__buf_1 _14024_ (.A(_07392_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_2 _14025_ (.A0(\core.cpuregs[11][23] ),
    .A1(_07239_),
    .S(_07389_),
    .X(_07393_));
 sky130_fd_sc_hd__buf_1 _14026_ (.A(_07393_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_2 _14027_ (.A0(\core.cpuregs[11][24] ),
    .A1(_07241_),
    .S(_07389_),
    .X(_07394_));
 sky130_fd_sc_hd__buf_1 _14028_ (.A(_07394_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_2 _14029_ (.A0(\core.cpuregs[11][25] ),
    .A1(_07243_),
    .S(_07389_),
    .X(_07395_));
 sky130_fd_sc_hd__buf_1 _14030_ (.A(_07395_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_2 _14031_ (.A0(\core.cpuregs[11][26] ),
    .A1(_07245_),
    .S(_07389_),
    .X(_07396_));
 sky130_fd_sc_hd__buf_1 _14032_ (.A(_07396_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_2 _14033_ (.A0(\core.cpuregs[11][27] ),
    .A1(_07247_),
    .S(_07389_),
    .X(_07397_));
 sky130_fd_sc_hd__buf_1 _14034_ (.A(_07397_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_2 _14035_ (.A0(\core.cpuregs[11][28] ),
    .A1(_07249_),
    .S(_07389_),
    .X(_07398_));
 sky130_fd_sc_hd__buf_1 _14036_ (.A(_07398_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_2 _14037_ (.A0(\core.cpuregs[11][29] ),
    .A1(_07251_),
    .S(_07389_),
    .X(_07399_));
 sky130_fd_sc_hd__buf_1 _14038_ (.A(_07399_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_2 _14039_ (.A0(\core.cpuregs[11][30] ),
    .A1(_07253_),
    .S(_07366_),
    .X(_07400_));
 sky130_fd_sc_hd__buf_1 _14040_ (.A(_07400_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_2 _14041_ (.A0(\core.cpuregs[11][31] ),
    .A1(_07255_),
    .S(_07366_),
    .X(_07401_));
 sky130_fd_sc_hd__buf_1 _14042_ (.A(_07401_),
    .X(_01022_));
 sky130_fd_sc_hd__or2_2 _14043_ (.A(_05464_),
    .B(_07365_),
    .X(_07402_));
 sky130_fd_sc_hd__buf_1 _14044_ (.A(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__mux2_2 _14045_ (.A0(_05460_),
    .A1(\core.cpuregs[10][0] ),
    .S(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__buf_1 _14046_ (.A(_07404_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_2 _14047_ (.A0(_05468_),
    .A1(\core.cpuregs[10][1] ),
    .S(_07403_),
    .X(_07405_));
 sky130_fd_sc_hd__buf_1 _14048_ (.A(_07405_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_2 _14049_ (.A0(_05470_),
    .A1(\core.cpuregs[10][2] ),
    .S(_07403_),
    .X(_07406_));
 sky130_fd_sc_hd__buf_1 _14050_ (.A(_07406_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_2 _14051_ (.A0(_05472_),
    .A1(\core.cpuregs[10][3] ),
    .S(_07403_),
    .X(_07407_));
 sky130_fd_sc_hd__buf_1 _14052_ (.A(_07407_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_2 _14053_ (.A0(_05474_),
    .A1(\core.cpuregs[10][4] ),
    .S(_07403_),
    .X(_07408_));
 sky130_fd_sc_hd__buf_1 _14054_ (.A(_07408_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_2 _14055_ (.A0(_05476_),
    .A1(\core.cpuregs[10][5] ),
    .S(_07403_),
    .X(_07409_));
 sky130_fd_sc_hd__buf_1 _14056_ (.A(_07409_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_2 _14057_ (.A0(_05478_),
    .A1(\core.cpuregs[10][6] ),
    .S(_07403_),
    .X(_07410_));
 sky130_fd_sc_hd__buf_1 _14058_ (.A(_07410_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_2 _14059_ (.A0(_05480_),
    .A1(\core.cpuregs[10][7] ),
    .S(_07403_),
    .X(_07411_));
 sky130_fd_sc_hd__buf_1 _14060_ (.A(_07411_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_2 _14061_ (.A0(_05482_),
    .A1(\core.cpuregs[10][8] ),
    .S(_07403_),
    .X(_07412_));
 sky130_fd_sc_hd__buf_1 _14062_ (.A(_07412_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_2 _14063_ (.A0(_05484_),
    .A1(\core.cpuregs[10][9] ),
    .S(_07403_),
    .X(_07413_));
 sky130_fd_sc_hd__buf_1 _14064_ (.A(_07413_),
    .X(_01032_));
 sky130_fd_sc_hd__buf_1 _14065_ (.A(_07402_),
    .X(_07414_));
 sky130_fd_sc_hd__mux2_2 _14066_ (.A0(_05486_),
    .A1(\core.cpuregs[10][10] ),
    .S(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__buf_1 _14067_ (.A(_07415_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_2 _14068_ (.A0(_05489_),
    .A1(\core.cpuregs[10][11] ),
    .S(_07414_),
    .X(_07416_));
 sky130_fd_sc_hd__buf_1 _14069_ (.A(_07416_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_2 _14070_ (.A0(_05491_),
    .A1(\core.cpuregs[10][12] ),
    .S(_07414_),
    .X(_07417_));
 sky130_fd_sc_hd__buf_1 _14071_ (.A(_07417_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_2 _14072_ (.A0(_05493_),
    .A1(\core.cpuregs[10][13] ),
    .S(_07414_),
    .X(_07418_));
 sky130_fd_sc_hd__buf_1 _14073_ (.A(_07418_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_2 _14074_ (.A0(_05495_),
    .A1(\core.cpuregs[10][14] ),
    .S(_07414_),
    .X(_07419_));
 sky130_fd_sc_hd__buf_1 _14075_ (.A(_07419_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_2 _14076_ (.A0(_05497_),
    .A1(\core.cpuregs[10][15] ),
    .S(_07414_),
    .X(_07420_));
 sky130_fd_sc_hd__buf_1 _14077_ (.A(_07420_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_2 _14078_ (.A0(_05499_),
    .A1(\core.cpuregs[10][16] ),
    .S(_07414_),
    .X(_07421_));
 sky130_fd_sc_hd__buf_1 _14079_ (.A(_07421_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_2 _14080_ (.A0(_05501_),
    .A1(\core.cpuregs[10][17] ),
    .S(_07414_),
    .X(_07422_));
 sky130_fd_sc_hd__buf_1 _14081_ (.A(_07422_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_2 _14082_ (.A0(_05503_),
    .A1(\core.cpuregs[10][18] ),
    .S(_07414_),
    .X(_07423_));
 sky130_fd_sc_hd__buf_1 _14083_ (.A(_07423_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_2 _14084_ (.A0(_05505_),
    .A1(\core.cpuregs[10][19] ),
    .S(_07414_),
    .X(_07424_));
 sky130_fd_sc_hd__buf_1 _14085_ (.A(_07424_),
    .X(_01042_));
 sky130_fd_sc_hd__buf_1 _14086_ (.A(_07402_),
    .X(_07425_));
 sky130_fd_sc_hd__mux2_2 _14087_ (.A0(_05507_),
    .A1(\core.cpuregs[10][20] ),
    .S(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__buf_1 _14088_ (.A(_07426_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_2 _14089_ (.A0(_05510_),
    .A1(\core.cpuregs[10][21] ),
    .S(_07425_),
    .X(_07427_));
 sky130_fd_sc_hd__buf_1 _14090_ (.A(_07427_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_2 _14091_ (.A0(_05512_),
    .A1(\core.cpuregs[10][22] ),
    .S(_07425_),
    .X(_07428_));
 sky130_fd_sc_hd__buf_1 _14092_ (.A(_07428_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_2 _14093_ (.A0(_05514_),
    .A1(\core.cpuregs[10][23] ),
    .S(_07425_),
    .X(_07429_));
 sky130_fd_sc_hd__buf_1 _14094_ (.A(_07429_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_2 _14095_ (.A0(_05516_),
    .A1(\core.cpuregs[10][24] ),
    .S(_07425_),
    .X(_07430_));
 sky130_fd_sc_hd__buf_1 _14096_ (.A(_07430_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_2 _14097_ (.A0(_05518_),
    .A1(\core.cpuregs[10][25] ),
    .S(_07425_),
    .X(_07431_));
 sky130_fd_sc_hd__buf_1 _14098_ (.A(_07431_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_2 _14099_ (.A0(_05520_),
    .A1(\core.cpuregs[10][26] ),
    .S(_07425_),
    .X(_07432_));
 sky130_fd_sc_hd__buf_1 _14100_ (.A(_07432_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_2 _14101_ (.A0(_05522_),
    .A1(\core.cpuregs[10][27] ),
    .S(_07425_),
    .X(_07433_));
 sky130_fd_sc_hd__buf_1 _14102_ (.A(_07433_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_2 _14103_ (.A0(_05524_),
    .A1(\core.cpuregs[10][28] ),
    .S(_07425_),
    .X(_07434_));
 sky130_fd_sc_hd__buf_1 _14104_ (.A(_07434_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_2 _14105_ (.A0(_05526_),
    .A1(\core.cpuregs[10][29] ),
    .S(_07425_),
    .X(_07435_));
 sky130_fd_sc_hd__buf_1 _14106_ (.A(_07435_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_2 _14107_ (.A0(_05528_),
    .A1(\core.cpuregs[10][30] ),
    .S(_07402_),
    .X(_07436_));
 sky130_fd_sc_hd__buf_1 _14108_ (.A(_07436_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_2 _14109_ (.A0(_05530_),
    .A1(\core.cpuregs[10][31] ),
    .S(_07402_),
    .X(_07437_));
 sky130_fd_sc_hd__buf_1 _14110_ (.A(_07437_),
    .X(_01054_));
 sky130_fd_sc_hd__buf_1 _14111_ (.A(\core.cpuregs[0][0] ),
    .X(_07438_));
 sky130_fd_sc_hd__buf_1 _14112_ (.A(_07438_),
    .X(_01055_));
 sky130_fd_sc_hd__buf_1 _14113_ (.A(\core.cpuregs[0][1] ),
    .X(_07439_));
 sky130_fd_sc_hd__buf_1 _14114_ (.A(_07439_),
    .X(_01056_));
 sky130_fd_sc_hd__buf_1 _14115_ (.A(\core.cpuregs[0][2] ),
    .X(_07440_));
 sky130_fd_sc_hd__buf_1 _14116_ (.A(_07440_),
    .X(_01057_));
 sky130_fd_sc_hd__buf_1 _14117_ (.A(\core.cpuregs[0][3] ),
    .X(_07441_));
 sky130_fd_sc_hd__buf_1 _14118_ (.A(_07441_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_1 _14119_ (.A(\core.cpuregs[0][4] ),
    .X(_07442_));
 sky130_fd_sc_hd__buf_1 _14120_ (.A(_07442_),
    .X(_01059_));
 sky130_fd_sc_hd__buf_1 _14121_ (.A(\core.cpuregs[0][5] ),
    .X(_07443_));
 sky130_fd_sc_hd__buf_1 _14122_ (.A(_07443_),
    .X(_01060_));
 sky130_fd_sc_hd__buf_1 _14123_ (.A(\core.cpuregs[0][6] ),
    .X(_07444_));
 sky130_fd_sc_hd__buf_1 _14124_ (.A(_07444_),
    .X(_01061_));
 sky130_fd_sc_hd__buf_1 _14125_ (.A(\core.cpuregs[0][7] ),
    .X(_07445_));
 sky130_fd_sc_hd__buf_1 _14126_ (.A(_07445_),
    .X(_01062_));
 sky130_fd_sc_hd__buf_1 _14127_ (.A(\core.cpuregs[0][8] ),
    .X(_07446_));
 sky130_fd_sc_hd__buf_1 _14128_ (.A(_07446_),
    .X(_01063_));
 sky130_fd_sc_hd__buf_1 _14129_ (.A(\core.cpuregs[0][9] ),
    .X(_07447_));
 sky130_fd_sc_hd__buf_1 _14130_ (.A(_07447_),
    .X(_01064_));
 sky130_fd_sc_hd__buf_1 _14131_ (.A(\core.cpuregs[0][10] ),
    .X(_07448_));
 sky130_fd_sc_hd__buf_1 _14132_ (.A(_07448_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_1 _14133_ (.A(\core.cpuregs[0][11] ),
    .X(_07449_));
 sky130_fd_sc_hd__buf_1 _14134_ (.A(_07449_),
    .X(_01066_));
 sky130_fd_sc_hd__buf_1 _14135_ (.A(\core.cpuregs[0][12] ),
    .X(_07450_));
 sky130_fd_sc_hd__buf_1 _14136_ (.A(_07450_),
    .X(_01067_));
 sky130_fd_sc_hd__buf_1 _14137_ (.A(\core.cpuregs[0][13] ),
    .X(_07451_));
 sky130_fd_sc_hd__buf_1 _14138_ (.A(_07451_),
    .X(_01068_));
 sky130_fd_sc_hd__buf_1 _14139_ (.A(\core.cpuregs[0][14] ),
    .X(_07452_));
 sky130_fd_sc_hd__buf_1 _14140_ (.A(_07452_),
    .X(_01069_));
 sky130_fd_sc_hd__buf_1 _14141_ (.A(\core.cpuregs[0][15] ),
    .X(_07453_));
 sky130_fd_sc_hd__buf_1 _14142_ (.A(_07453_),
    .X(_01070_));
 sky130_fd_sc_hd__buf_1 _14143_ (.A(\core.cpuregs[0][16] ),
    .X(_07454_));
 sky130_fd_sc_hd__buf_1 _14144_ (.A(_07454_),
    .X(_01071_));
 sky130_fd_sc_hd__buf_1 _14145_ (.A(\core.cpuregs[0][17] ),
    .X(_07455_));
 sky130_fd_sc_hd__buf_1 _14146_ (.A(_07455_),
    .X(_01072_));
 sky130_fd_sc_hd__buf_1 _14147_ (.A(\core.cpuregs[0][18] ),
    .X(_07456_));
 sky130_fd_sc_hd__buf_1 _14148_ (.A(_07456_),
    .X(_01073_));
 sky130_fd_sc_hd__buf_1 _14149_ (.A(\core.cpuregs[0][19] ),
    .X(_07457_));
 sky130_fd_sc_hd__buf_1 _14150_ (.A(_07457_),
    .X(_01074_));
 sky130_fd_sc_hd__buf_1 _14151_ (.A(\core.cpuregs[0][20] ),
    .X(_07458_));
 sky130_fd_sc_hd__buf_1 _14152_ (.A(_07458_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_1 _14153_ (.A(\core.cpuregs[0][21] ),
    .X(_07459_));
 sky130_fd_sc_hd__buf_1 _14154_ (.A(_07459_),
    .X(_01076_));
 sky130_fd_sc_hd__buf_1 _14155_ (.A(\core.cpuregs[0][22] ),
    .X(_07460_));
 sky130_fd_sc_hd__buf_1 _14156_ (.A(_07460_),
    .X(_01077_));
 sky130_fd_sc_hd__buf_1 _14157_ (.A(\core.cpuregs[0][23] ),
    .X(_07461_));
 sky130_fd_sc_hd__buf_1 _14158_ (.A(_07461_),
    .X(_01078_));
 sky130_fd_sc_hd__buf_1 _14159_ (.A(\core.cpuregs[0][24] ),
    .X(_07462_));
 sky130_fd_sc_hd__buf_1 _14160_ (.A(_07462_),
    .X(_01079_));
 sky130_fd_sc_hd__buf_1 _14161_ (.A(\core.cpuregs[0][25] ),
    .X(_07463_));
 sky130_fd_sc_hd__buf_1 _14162_ (.A(_07463_),
    .X(_01080_));
 sky130_fd_sc_hd__buf_1 _14163_ (.A(\core.cpuregs[0][26] ),
    .X(_07464_));
 sky130_fd_sc_hd__buf_1 _14164_ (.A(_07464_),
    .X(_01081_));
 sky130_fd_sc_hd__buf_1 _14165_ (.A(\core.cpuregs[0][27] ),
    .X(_07465_));
 sky130_fd_sc_hd__buf_1 _14166_ (.A(_07465_),
    .X(_01082_));
 sky130_fd_sc_hd__buf_1 _14167_ (.A(\core.cpuregs[0][28] ),
    .X(_07466_));
 sky130_fd_sc_hd__buf_1 _14168_ (.A(_07466_),
    .X(_01083_));
 sky130_fd_sc_hd__buf_1 _14169_ (.A(\core.cpuregs[0][29] ),
    .X(_07467_));
 sky130_fd_sc_hd__buf_1 _14170_ (.A(_07467_),
    .X(_01084_));
 sky130_fd_sc_hd__buf_1 _14171_ (.A(\core.cpuregs[0][30] ),
    .X(_07468_));
 sky130_fd_sc_hd__buf_1 _14172_ (.A(_07468_),
    .X(_01085_));
 sky130_fd_sc_hd__buf_1 _14173_ (.A(\core.cpuregs[0][31] ),
    .X(_07469_));
 sky130_fd_sc_hd__buf_1 _14174_ (.A(_07469_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_2 _14175_ (.A(_05766_),
    .B(_07365_),
    .X(_07470_));
 sky130_fd_sc_hd__buf_1 _14176_ (.A(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__mux2_2 _14177_ (.A0(_05460_),
    .A1(\core.cpuregs[8][0] ),
    .S(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__buf_1 _14178_ (.A(_07472_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_2 _14179_ (.A0(_05468_),
    .A1(\core.cpuregs[8][1] ),
    .S(_07471_),
    .X(_07473_));
 sky130_fd_sc_hd__buf_1 _14180_ (.A(_07473_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_2 _14181_ (.A0(_05470_),
    .A1(\core.cpuregs[8][2] ),
    .S(_07471_),
    .X(_07474_));
 sky130_fd_sc_hd__buf_1 _14182_ (.A(_07474_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_2 _14183_ (.A0(_05472_),
    .A1(\core.cpuregs[8][3] ),
    .S(_07471_),
    .X(_07475_));
 sky130_fd_sc_hd__buf_1 _14184_ (.A(_07475_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_2 _14185_ (.A0(_05474_),
    .A1(\core.cpuregs[8][4] ),
    .S(_07471_),
    .X(_07476_));
 sky130_fd_sc_hd__buf_1 _14186_ (.A(_07476_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_2 _14187_ (.A0(_05476_),
    .A1(\core.cpuregs[8][5] ),
    .S(_07471_),
    .X(_07477_));
 sky130_fd_sc_hd__buf_1 _14188_ (.A(_07477_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_2 _14189_ (.A0(_05478_),
    .A1(\core.cpuregs[8][6] ),
    .S(_07471_),
    .X(_07478_));
 sky130_fd_sc_hd__buf_1 _14190_ (.A(_07478_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_2 _14191_ (.A0(_05480_),
    .A1(\core.cpuregs[8][7] ),
    .S(_07471_),
    .X(_07479_));
 sky130_fd_sc_hd__buf_1 _14192_ (.A(_07479_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_2 _14193_ (.A0(_05482_),
    .A1(\core.cpuregs[8][8] ),
    .S(_07471_),
    .X(_07480_));
 sky130_fd_sc_hd__buf_1 _14194_ (.A(_07480_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_2 _14195_ (.A0(_05484_),
    .A1(\core.cpuregs[8][9] ),
    .S(_07471_),
    .X(_07481_));
 sky130_fd_sc_hd__buf_1 _14196_ (.A(_07481_),
    .X(_01096_));
 sky130_fd_sc_hd__buf_1 _14197_ (.A(_07470_),
    .X(_07482_));
 sky130_fd_sc_hd__mux2_2 _14198_ (.A0(_05486_),
    .A1(\core.cpuregs[8][10] ),
    .S(_07482_),
    .X(_07483_));
 sky130_fd_sc_hd__buf_1 _14199_ (.A(_07483_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_2 _14200_ (.A0(_05489_),
    .A1(\core.cpuregs[8][11] ),
    .S(_07482_),
    .X(_07484_));
 sky130_fd_sc_hd__buf_1 _14201_ (.A(_07484_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_2 _14202_ (.A0(_05491_),
    .A1(\core.cpuregs[8][12] ),
    .S(_07482_),
    .X(_07485_));
 sky130_fd_sc_hd__buf_1 _14203_ (.A(_07485_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_2 _14204_ (.A0(_05493_),
    .A1(\core.cpuregs[8][13] ),
    .S(_07482_),
    .X(_07486_));
 sky130_fd_sc_hd__buf_1 _14205_ (.A(_07486_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_2 _14206_ (.A0(_05495_),
    .A1(\core.cpuregs[8][14] ),
    .S(_07482_),
    .X(_07487_));
 sky130_fd_sc_hd__buf_1 _14207_ (.A(_07487_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_2 _14208_ (.A0(_05497_),
    .A1(\core.cpuregs[8][15] ),
    .S(_07482_),
    .X(_07488_));
 sky130_fd_sc_hd__buf_1 _14209_ (.A(_07488_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_2 _14210_ (.A0(_05499_),
    .A1(\core.cpuregs[8][16] ),
    .S(_07482_),
    .X(_07489_));
 sky130_fd_sc_hd__buf_1 _14211_ (.A(_07489_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_2 _14212_ (.A0(_05501_),
    .A1(\core.cpuregs[8][17] ),
    .S(_07482_),
    .X(_07490_));
 sky130_fd_sc_hd__buf_1 _14213_ (.A(_07490_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_2 _14214_ (.A0(_05503_),
    .A1(\core.cpuregs[8][18] ),
    .S(_07482_),
    .X(_07491_));
 sky130_fd_sc_hd__buf_1 _14215_ (.A(_07491_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_2 _14216_ (.A0(_05505_),
    .A1(\core.cpuregs[8][19] ),
    .S(_07482_),
    .X(_07492_));
 sky130_fd_sc_hd__buf_1 _14217_ (.A(_07492_),
    .X(_01106_));
 sky130_fd_sc_hd__buf_1 _14218_ (.A(_07470_),
    .X(_07493_));
 sky130_fd_sc_hd__mux2_2 _14219_ (.A0(_05507_),
    .A1(\core.cpuregs[8][20] ),
    .S(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__buf_1 _14220_ (.A(_07494_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_2 _14221_ (.A0(_05510_),
    .A1(\core.cpuregs[8][21] ),
    .S(_07493_),
    .X(_07495_));
 sky130_fd_sc_hd__buf_1 _14222_ (.A(_07495_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_2 _14223_ (.A0(_05512_),
    .A1(\core.cpuregs[8][22] ),
    .S(_07493_),
    .X(_07496_));
 sky130_fd_sc_hd__buf_1 _14224_ (.A(_07496_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_2 _14225_ (.A0(_05514_),
    .A1(\core.cpuregs[8][23] ),
    .S(_07493_),
    .X(_07497_));
 sky130_fd_sc_hd__buf_1 _14226_ (.A(_07497_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_2 _14227_ (.A0(_05516_),
    .A1(\core.cpuregs[8][24] ),
    .S(_07493_),
    .X(_07498_));
 sky130_fd_sc_hd__buf_1 _14228_ (.A(_07498_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_2 _14229_ (.A0(_05518_),
    .A1(\core.cpuregs[8][25] ),
    .S(_07493_),
    .X(_07499_));
 sky130_fd_sc_hd__buf_1 _14230_ (.A(_07499_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_2 _14231_ (.A0(_05520_),
    .A1(\core.cpuregs[8][26] ),
    .S(_07493_),
    .X(_07500_));
 sky130_fd_sc_hd__buf_1 _14232_ (.A(_07500_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_2 _14233_ (.A0(_05522_),
    .A1(\core.cpuregs[8][27] ),
    .S(_07493_),
    .X(_07501_));
 sky130_fd_sc_hd__buf_1 _14234_ (.A(_07501_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_2 _14235_ (.A0(_05524_),
    .A1(\core.cpuregs[8][28] ),
    .S(_07493_),
    .X(_07502_));
 sky130_fd_sc_hd__buf_1 _14236_ (.A(_07502_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_2 _14237_ (.A0(_05526_),
    .A1(\core.cpuregs[8][29] ),
    .S(_07493_),
    .X(_07503_));
 sky130_fd_sc_hd__buf_1 _14238_ (.A(_07503_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_2 _14239_ (.A0(_05528_),
    .A1(\core.cpuregs[8][30] ),
    .S(_07470_),
    .X(_07504_));
 sky130_fd_sc_hd__buf_1 _14240_ (.A(_07504_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_2 _14241_ (.A0(_05530_),
    .A1(\core.cpuregs[8][31] ),
    .S(_07470_),
    .X(_07505_));
 sky130_fd_sc_hd__buf_1 _14242_ (.A(_07505_),
    .X(_01118_));
 sky130_fd_sc_hd__or3b_2 _14243_ (.A(\core.latched_rd[4] ),
    .B(\core.latched_rd[3] ),
    .C_N(\core.latched_rd[2] ),
    .X(_07506_));
 sky130_fd_sc_hd__nor2_2 _14244_ (.A(_05286_),
    .B(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__buf_1 _14245_ (.A(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__mux2_2 _14246_ (.A0(\core.cpuregs[7][0] ),
    .A1(_07188_),
    .S(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__buf_1 _14247_ (.A(_07509_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_2 _14248_ (.A0(\core.cpuregs[7][1] ),
    .A1(_07193_),
    .S(_07508_),
    .X(_07510_));
 sky130_fd_sc_hd__buf_1 _14249_ (.A(_07510_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_2 _14250_ (.A0(\core.cpuregs[7][2] ),
    .A1(_07195_),
    .S(_07508_),
    .X(_07511_));
 sky130_fd_sc_hd__buf_1 _14251_ (.A(_07511_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_2 _14252_ (.A0(\core.cpuregs[7][3] ),
    .A1(_07197_),
    .S(_07508_),
    .X(_07512_));
 sky130_fd_sc_hd__buf_1 _14253_ (.A(_07512_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_2 _14254_ (.A0(\core.cpuregs[7][4] ),
    .A1(_07199_),
    .S(_07508_),
    .X(_07513_));
 sky130_fd_sc_hd__buf_1 _14255_ (.A(_07513_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_2 _14256_ (.A0(\core.cpuregs[7][5] ),
    .A1(_07201_),
    .S(_07508_),
    .X(_07514_));
 sky130_fd_sc_hd__buf_1 _14257_ (.A(_07514_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_2 _14258_ (.A0(\core.cpuregs[7][6] ),
    .A1(_07203_),
    .S(_07508_),
    .X(_07515_));
 sky130_fd_sc_hd__buf_1 _14259_ (.A(_07515_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_2 _14260_ (.A0(\core.cpuregs[7][7] ),
    .A1(_07205_),
    .S(_07508_),
    .X(_07516_));
 sky130_fd_sc_hd__buf_1 _14261_ (.A(_07516_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_2 _14262_ (.A0(\core.cpuregs[7][8] ),
    .A1(_07207_),
    .S(_07508_),
    .X(_07517_));
 sky130_fd_sc_hd__buf_1 _14263_ (.A(_07517_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_2 _14264_ (.A0(\core.cpuregs[7][9] ),
    .A1(_07209_),
    .S(_07508_),
    .X(_07518_));
 sky130_fd_sc_hd__buf_1 _14265_ (.A(_07518_),
    .X(_01128_));
 sky130_fd_sc_hd__buf_1 _14266_ (.A(_07507_),
    .X(_07519_));
 sky130_fd_sc_hd__mux2_2 _14267_ (.A0(\core.cpuregs[7][10] ),
    .A1(_07211_),
    .S(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__buf_1 _14268_ (.A(_07520_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_2 _14269_ (.A0(\core.cpuregs[7][11] ),
    .A1(_07214_),
    .S(_07519_),
    .X(_07521_));
 sky130_fd_sc_hd__buf_1 _14270_ (.A(_07521_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_2 _14271_ (.A0(\core.cpuregs[7][12] ),
    .A1(_07216_),
    .S(_07519_),
    .X(_07522_));
 sky130_fd_sc_hd__buf_1 _14272_ (.A(_07522_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_2 _14273_ (.A0(\core.cpuregs[7][13] ),
    .A1(_07218_),
    .S(_07519_),
    .X(_07523_));
 sky130_fd_sc_hd__buf_1 _14274_ (.A(_07523_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_2 _14275_ (.A0(\core.cpuregs[7][14] ),
    .A1(_07220_),
    .S(_07519_),
    .X(_07524_));
 sky130_fd_sc_hd__buf_1 _14276_ (.A(_07524_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_2 _14277_ (.A0(\core.cpuregs[7][15] ),
    .A1(_07222_),
    .S(_07519_),
    .X(_07525_));
 sky130_fd_sc_hd__buf_1 _14278_ (.A(_07525_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_2 _14279_ (.A0(\core.cpuregs[7][16] ),
    .A1(_07224_),
    .S(_07519_),
    .X(_07526_));
 sky130_fd_sc_hd__buf_1 _14280_ (.A(_07526_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_2 _14281_ (.A0(\core.cpuregs[7][17] ),
    .A1(_07226_),
    .S(_07519_),
    .X(_07527_));
 sky130_fd_sc_hd__buf_1 _14282_ (.A(_07527_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_2 _14283_ (.A0(\core.cpuregs[7][18] ),
    .A1(_07228_),
    .S(_07519_),
    .X(_07528_));
 sky130_fd_sc_hd__buf_1 _14284_ (.A(_07528_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_2 _14285_ (.A0(\core.cpuregs[7][19] ),
    .A1(_07230_),
    .S(_07519_),
    .X(_07529_));
 sky130_fd_sc_hd__buf_1 _14286_ (.A(_07529_),
    .X(_01138_));
 sky130_fd_sc_hd__buf_1 _14287_ (.A(_07507_),
    .X(_07530_));
 sky130_fd_sc_hd__mux2_2 _14288_ (.A0(\core.cpuregs[7][20] ),
    .A1(_07232_),
    .S(_07530_),
    .X(_07531_));
 sky130_fd_sc_hd__buf_1 _14289_ (.A(_07531_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_2 _14290_ (.A0(\core.cpuregs[7][21] ),
    .A1(_07235_),
    .S(_07530_),
    .X(_07532_));
 sky130_fd_sc_hd__buf_1 _14291_ (.A(_07532_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_2 _14292_ (.A0(\core.cpuregs[7][22] ),
    .A1(_07237_),
    .S(_07530_),
    .X(_07533_));
 sky130_fd_sc_hd__buf_1 _14293_ (.A(_07533_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_2 _14294_ (.A0(\core.cpuregs[7][23] ),
    .A1(_07239_),
    .S(_07530_),
    .X(_07534_));
 sky130_fd_sc_hd__buf_1 _14295_ (.A(_07534_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_2 _14296_ (.A0(\core.cpuregs[7][24] ),
    .A1(_07241_),
    .S(_07530_),
    .X(_07535_));
 sky130_fd_sc_hd__buf_1 _14297_ (.A(_07535_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_2 _14298_ (.A0(\core.cpuregs[7][25] ),
    .A1(_07243_),
    .S(_07530_),
    .X(_07536_));
 sky130_fd_sc_hd__buf_1 _14299_ (.A(_07536_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_2 _14300_ (.A0(\core.cpuregs[7][26] ),
    .A1(_07245_),
    .S(_07530_),
    .X(_07537_));
 sky130_fd_sc_hd__buf_1 _14301_ (.A(_07537_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_2 _14302_ (.A0(\core.cpuregs[7][27] ),
    .A1(_07247_),
    .S(_07530_),
    .X(_07538_));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(_07538_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_2 _14304_ (.A0(\core.cpuregs[7][28] ),
    .A1(_07249_),
    .S(_07530_),
    .X(_07539_));
 sky130_fd_sc_hd__buf_1 _14305_ (.A(_07539_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_2 _14306_ (.A0(\core.cpuregs[7][29] ),
    .A1(_07251_),
    .S(_07530_),
    .X(_07540_));
 sky130_fd_sc_hd__buf_1 _14307_ (.A(_07540_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_2 _14308_ (.A0(\core.cpuregs[7][30] ),
    .A1(_07253_),
    .S(_07507_),
    .X(_07541_));
 sky130_fd_sc_hd__buf_1 _14309_ (.A(_07541_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_2 _14310_ (.A0(\core.cpuregs[7][31] ),
    .A1(_07255_),
    .S(_07507_),
    .X(_07542_));
 sky130_fd_sc_hd__buf_1 _14311_ (.A(_07542_),
    .X(_01150_));
 sky130_fd_sc_hd__or2_2 _14312_ (.A(_05464_),
    .B(_07506_),
    .X(_07543_));
 sky130_fd_sc_hd__buf_1 _14313_ (.A(_07543_),
    .X(_07544_));
 sky130_fd_sc_hd__mux2_2 _14314_ (.A0(_05284_),
    .A1(\core.cpuregs[6][0] ),
    .S(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__buf_1 _14315_ (.A(_07545_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_2 _14316_ (.A0(_05292_),
    .A1(\core.cpuregs[6][1] ),
    .S(_07544_),
    .X(_07546_));
 sky130_fd_sc_hd__buf_1 _14317_ (.A(_07546_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_2 _14318_ (.A0(_05297_),
    .A1(\core.cpuregs[6][2] ),
    .S(_07544_),
    .X(_07547_));
 sky130_fd_sc_hd__buf_1 _14319_ (.A(_07547_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_2 _14320_ (.A0(_05304_),
    .A1(\core.cpuregs[6][3] ),
    .S(_07544_),
    .X(_01575_));
 sky130_fd_sc_hd__buf_1 _14321_ (.A(_01575_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_2 _14322_ (.A0(_05310_),
    .A1(\core.cpuregs[6][4] ),
    .S(_07544_),
    .X(_01576_));
 sky130_fd_sc_hd__buf_1 _14323_ (.A(_01576_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_2 _14324_ (.A0(_05315_),
    .A1(\core.cpuregs[6][5] ),
    .S(_07544_),
    .X(_01577_));
 sky130_fd_sc_hd__buf_1 _14325_ (.A(_01577_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_2 _14326_ (.A0(_05320_),
    .A1(\core.cpuregs[6][6] ),
    .S(_07544_),
    .X(_01578_));
 sky130_fd_sc_hd__buf_1 _14327_ (.A(_01578_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_2 _14328_ (.A0(_05326_),
    .A1(\core.cpuregs[6][7] ),
    .S(_07544_),
    .X(_01579_));
 sky130_fd_sc_hd__buf_1 _14329_ (.A(_01579_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_2 _14330_ (.A0(_05332_),
    .A1(\core.cpuregs[6][8] ),
    .S(_07544_),
    .X(_01580_));
 sky130_fd_sc_hd__buf_1 _14331_ (.A(_01580_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_2 _14332_ (.A0(_05337_),
    .A1(\core.cpuregs[6][9] ),
    .S(_07544_),
    .X(_01581_));
 sky130_fd_sc_hd__buf_1 _14333_ (.A(_01581_),
    .X(_01160_));
 sky130_fd_sc_hd__buf_1 _14334_ (.A(_07543_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_2 _14335_ (.A0(_05343_),
    .A1(\core.cpuregs[6][10] ),
    .S(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__buf_1 _14336_ (.A(_01583_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_2 _14337_ (.A0(_05349_),
    .A1(\core.cpuregs[6][11] ),
    .S(_01582_),
    .X(_01584_));
 sky130_fd_sc_hd__buf_1 _14338_ (.A(_01584_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_2 _14339_ (.A0(_05355_),
    .A1(\core.cpuregs[6][12] ),
    .S(_01582_),
    .X(_01585_));
 sky130_fd_sc_hd__buf_1 _14340_ (.A(_01585_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_2 _14341_ (.A0(_05360_),
    .A1(\core.cpuregs[6][13] ),
    .S(_01582_),
    .X(_01586_));
 sky130_fd_sc_hd__buf_1 _14342_ (.A(_01586_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_2 _14343_ (.A0(_05367_),
    .A1(\core.cpuregs[6][14] ),
    .S(_01582_),
    .X(_01587_));
 sky130_fd_sc_hd__buf_1 _14344_ (.A(_01587_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_2 _14345_ (.A0(_05372_),
    .A1(\core.cpuregs[6][15] ),
    .S(_01582_),
    .X(_01588_));
 sky130_fd_sc_hd__buf_1 _14346_ (.A(_01588_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_2 _14347_ (.A0(_05377_),
    .A1(\core.cpuregs[6][16] ),
    .S(_01582_),
    .X(_01589_));
 sky130_fd_sc_hd__buf_1 _14348_ (.A(_01589_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_2 _14349_ (.A0(_05383_),
    .A1(\core.cpuregs[6][17] ),
    .S(_01582_),
    .X(_01590_));
 sky130_fd_sc_hd__buf_1 _14350_ (.A(_01590_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_2 _14351_ (.A0(_05388_),
    .A1(\core.cpuregs[6][18] ),
    .S(_01582_),
    .X(_01591_));
 sky130_fd_sc_hd__buf_1 _14352_ (.A(_01591_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_2 _14353_ (.A0(_05393_),
    .A1(\core.cpuregs[6][19] ),
    .S(_01582_),
    .X(_01592_));
 sky130_fd_sc_hd__buf_1 _14354_ (.A(_01592_),
    .X(_01170_));
 sky130_fd_sc_hd__buf_1 _14355_ (.A(_07543_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_2 _14356_ (.A0(_05399_),
    .A1(\core.cpuregs[6][20] ),
    .S(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_1 _14357_ (.A(_01594_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_2 _14358_ (.A0(_05405_),
    .A1(\core.cpuregs[6][21] ),
    .S(_01593_),
    .X(_01595_));
 sky130_fd_sc_hd__buf_1 _14359_ (.A(_01595_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_2 _14360_ (.A0(_05410_),
    .A1(\core.cpuregs[6][22] ),
    .S(_01593_),
    .X(_01596_));
 sky130_fd_sc_hd__buf_1 _14361_ (.A(_01596_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_2 _14362_ (.A0(_05416_),
    .A1(\core.cpuregs[6][23] ),
    .S(_01593_),
    .X(_01597_));
 sky130_fd_sc_hd__buf_1 _14363_ (.A(_01597_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_2 _14364_ (.A0(_05421_),
    .A1(\core.cpuregs[6][24] ),
    .S(_01593_),
    .X(_01598_));
 sky130_fd_sc_hd__buf_1 _14365_ (.A(_01598_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_2 _14366_ (.A0(_05426_),
    .A1(\core.cpuregs[6][25] ),
    .S(_01593_),
    .X(_01599_));
 sky130_fd_sc_hd__buf_1 _14367_ (.A(_01599_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_2 _14368_ (.A0(_05432_),
    .A1(\core.cpuregs[6][26] ),
    .S(_01593_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_1 _14369_ (.A(_01600_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_2 _14370_ (.A0(_05437_),
    .A1(\core.cpuregs[6][27] ),
    .S(_01593_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_1 _14371_ (.A(_01601_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_2 _14372_ (.A0(_05442_),
    .A1(\core.cpuregs[6][28] ),
    .S(_01593_),
    .X(_01602_));
 sky130_fd_sc_hd__buf_1 _14373_ (.A(_01602_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_2 _14374_ (.A0(_05448_),
    .A1(\core.cpuregs[6][29] ),
    .S(_01593_),
    .X(_01603_));
 sky130_fd_sc_hd__buf_1 _14375_ (.A(_01603_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_2 _14376_ (.A0(_05453_),
    .A1(\core.cpuregs[6][30] ),
    .S(_07543_),
    .X(_01604_));
 sky130_fd_sc_hd__buf_1 _14377_ (.A(_01604_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_2 _14378_ (.A0(_05458_),
    .A1(\core.cpuregs[6][31] ),
    .S(_07543_),
    .X(_01605_));
 sky130_fd_sc_hd__buf_1 _14379_ (.A(_01605_),
    .X(_01182_));
 sky130_fd_sc_hd__or2_2 _14380_ (.A(_05837_),
    .B(_07506_),
    .X(_01606_));
 sky130_fd_sc_hd__buf_1 _14381_ (.A(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_2 _14382_ (.A0(_05284_),
    .A1(\core.cpuregs[5][0] ),
    .S(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_1 _14383_ (.A(_01608_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_2 _14384_ (.A0(_05292_),
    .A1(\core.cpuregs[5][1] ),
    .S(_01607_),
    .X(_01609_));
 sky130_fd_sc_hd__buf_1 _14385_ (.A(_01609_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_2 _14386_ (.A0(_05297_),
    .A1(\core.cpuregs[5][2] ),
    .S(_01607_),
    .X(_01610_));
 sky130_fd_sc_hd__buf_1 _14387_ (.A(_01610_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_2 _14388_ (.A0(_05304_),
    .A1(\core.cpuregs[5][3] ),
    .S(_01607_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_1 _14389_ (.A(_01611_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_2 _14390_ (.A0(_05310_),
    .A1(\core.cpuregs[5][4] ),
    .S(_01607_),
    .X(_01612_));
 sky130_fd_sc_hd__buf_1 _14391_ (.A(_01612_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_2 _14392_ (.A0(_05315_),
    .A1(\core.cpuregs[5][5] ),
    .S(_01607_),
    .X(_01613_));
 sky130_fd_sc_hd__buf_1 _14393_ (.A(_01613_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_2 _14394_ (.A0(_05320_),
    .A1(\core.cpuregs[5][6] ),
    .S(_01607_),
    .X(_01614_));
 sky130_fd_sc_hd__buf_1 _14395_ (.A(_01614_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_2 _14396_ (.A0(_05326_),
    .A1(\core.cpuregs[5][7] ),
    .S(_01607_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_1 _14397_ (.A(_01615_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_2 _14398_ (.A0(_05332_),
    .A1(\core.cpuregs[5][8] ),
    .S(_01607_),
    .X(_01616_));
 sky130_fd_sc_hd__buf_1 _14399_ (.A(_01616_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_2 _14400_ (.A0(_05337_),
    .A1(\core.cpuregs[5][9] ),
    .S(_01607_),
    .X(_01617_));
 sky130_fd_sc_hd__buf_1 _14401_ (.A(_01617_),
    .X(_01192_));
 sky130_fd_sc_hd__buf_1 _14402_ (.A(_01606_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_2 _14403_ (.A0(_05343_),
    .A1(\core.cpuregs[5][10] ),
    .S(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__buf_1 _14404_ (.A(_01619_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_2 _14405_ (.A0(_05349_),
    .A1(\core.cpuregs[5][11] ),
    .S(_01618_),
    .X(_01620_));
 sky130_fd_sc_hd__buf_1 _14406_ (.A(_01620_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_2 _14407_ (.A0(_05355_),
    .A1(\core.cpuregs[5][12] ),
    .S(_01618_),
    .X(_01621_));
 sky130_fd_sc_hd__buf_1 _14408_ (.A(_01621_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_2 _14409_ (.A0(_05360_),
    .A1(\core.cpuregs[5][13] ),
    .S(_01618_),
    .X(_01622_));
 sky130_fd_sc_hd__buf_1 _14410_ (.A(_01622_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_2 _14411_ (.A0(_05367_),
    .A1(\core.cpuregs[5][14] ),
    .S(_01618_),
    .X(_01623_));
 sky130_fd_sc_hd__buf_1 _14412_ (.A(_01623_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_2 _14413_ (.A0(_05372_),
    .A1(\core.cpuregs[5][15] ),
    .S(_01618_),
    .X(_01624_));
 sky130_fd_sc_hd__buf_1 _14414_ (.A(_01624_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_2 _14415_ (.A0(_05377_),
    .A1(\core.cpuregs[5][16] ),
    .S(_01618_),
    .X(_01625_));
 sky130_fd_sc_hd__buf_1 _14416_ (.A(_01625_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_2 _14417_ (.A0(_05383_),
    .A1(\core.cpuregs[5][17] ),
    .S(_01618_),
    .X(_01626_));
 sky130_fd_sc_hd__buf_1 _14418_ (.A(_01626_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_2 _14419_ (.A0(_05388_),
    .A1(\core.cpuregs[5][18] ),
    .S(_01618_),
    .X(_01627_));
 sky130_fd_sc_hd__buf_1 _14420_ (.A(_01627_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_2 _14421_ (.A0(_05393_),
    .A1(\core.cpuregs[5][19] ),
    .S(_01618_),
    .X(_01628_));
 sky130_fd_sc_hd__buf_1 _14422_ (.A(_01628_),
    .X(_01202_));
 sky130_fd_sc_hd__buf_1 _14423_ (.A(_01606_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_2 _14424_ (.A0(_05399_),
    .A1(\core.cpuregs[5][20] ),
    .S(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__buf_1 _14425_ (.A(_01630_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_2 _14426_ (.A0(_05405_),
    .A1(\core.cpuregs[5][21] ),
    .S(_01629_),
    .X(_01631_));
 sky130_fd_sc_hd__buf_1 _14427_ (.A(_01631_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_2 _14428_ (.A0(_05410_),
    .A1(\core.cpuregs[5][22] ),
    .S(_01629_),
    .X(_01632_));
 sky130_fd_sc_hd__buf_1 _14429_ (.A(_01632_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_2 _14430_ (.A0(_05416_),
    .A1(\core.cpuregs[5][23] ),
    .S(_01629_),
    .X(_01633_));
 sky130_fd_sc_hd__buf_1 _14431_ (.A(_01633_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_2 _14432_ (.A0(_05421_),
    .A1(\core.cpuregs[5][24] ),
    .S(_01629_),
    .X(_01634_));
 sky130_fd_sc_hd__buf_1 _14433_ (.A(_01634_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_2 _14434_ (.A0(_05426_),
    .A1(\core.cpuregs[5][25] ),
    .S(_01629_),
    .X(_01635_));
 sky130_fd_sc_hd__buf_1 _14435_ (.A(_01635_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_2 _14436_ (.A0(_05432_),
    .A1(\core.cpuregs[5][26] ),
    .S(_01629_),
    .X(_01636_));
 sky130_fd_sc_hd__buf_1 _14437_ (.A(_01636_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_2 _14438_ (.A0(_05437_),
    .A1(\core.cpuregs[5][27] ),
    .S(_01629_),
    .X(_01637_));
 sky130_fd_sc_hd__buf_1 _14439_ (.A(_01637_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_2 _14440_ (.A0(_05442_),
    .A1(\core.cpuregs[5][28] ),
    .S(_01629_),
    .X(_01638_));
 sky130_fd_sc_hd__buf_1 _14441_ (.A(_01638_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_2 _14442_ (.A0(_05448_),
    .A1(\core.cpuregs[5][29] ),
    .S(_01629_),
    .X(_01639_));
 sky130_fd_sc_hd__buf_1 _14443_ (.A(_01639_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_2 _14444_ (.A0(_05453_),
    .A1(\core.cpuregs[5][30] ),
    .S(_01606_),
    .X(_01640_));
 sky130_fd_sc_hd__buf_1 _14445_ (.A(_01640_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_2 _14446_ (.A0(_05458_),
    .A1(\core.cpuregs[5][31] ),
    .S(_01606_),
    .X(_01641_));
 sky130_fd_sc_hd__buf_1 _14447_ (.A(_01641_),
    .X(_01214_));
 sky130_fd_sc_hd__nor2_2 _14448_ (.A(_05766_),
    .B(_07506_),
    .Y(_01642_));
 sky130_fd_sc_hd__buf_1 _14449_ (.A(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_2 _14450_ (.A0(\core.cpuregs[4][0] ),
    .A1(_07188_),
    .S(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__buf_1 _14451_ (.A(_01644_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_2 _14452_ (.A0(\core.cpuregs[4][1] ),
    .A1(_07193_),
    .S(_01643_),
    .X(_01645_));
 sky130_fd_sc_hd__buf_1 _14453_ (.A(_01645_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_2 _14454_ (.A0(\core.cpuregs[4][2] ),
    .A1(_07195_),
    .S(_01643_),
    .X(_01646_));
 sky130_fd_sc_hd__buf_1 _14455_ (.A(_01646_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_2 _14456_ (.A0(\core.cpuregs[4][3] ),
    .A1(_07197_),
    .S(_01643_),
    .X(_01647_));
 sky130_fd_sc_hd__buf_1 _14457_ (.A(_01647_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_2 _14458_ (.A0(\core.cpuregs[4][4] ),
    .A1(_07199_),
    .S(_01643_),
    .X(_01648_));
 sky130_fd_sc_hd__buf_1 _14459_ (.A(_01648_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_2 _14460_ (.A0(\core.cpuregs[4][5] ),
    .A1(_07201_),
    .S(_01643_),
    .X(_01649_));
 sky130_fd_sc_hd__buf_1 _14461_ (.A(_01649_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_2 _14462_ (.A0(\core.cpuregs[4][6] ),
    .A1(_07203_),
    .S(_01643_),
    .X(_01650_));
 sky130_fd_sc_hd__buf_1 _14463_ (.A(_01650_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_2 _14464_ (.A0(\core.cpuregs[4][7] ),
    .A1(_07205_),
    .S(_01643_),
    .X(_01651_));
 sky130_fd_sc_hd__buf_1 _14465_ (.A(_01651_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_2 _14466_ (.A0(\core.cpuregs[4][8] ),
    .A1(_07207_),
    .S(_01643_),
    .X(_01652_));
 sky130_fd_sc_hd__buf_1 _14467_ (.A(_01652_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_2 _14468_ (.A0(\core.cpuregs[4][9] ),
    .A1(_07209_),
    .S(_01643_),
    .X(_01653_));
 sky130_fd_sc_hd__buf_1 _14469_ (.A(_01653_),
    .X(_01224_));
 sky130_fd_sc_hd__buf_1 _14470_ (.A(_01642_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_2 _14471_ (.A0(\core.cpuregs[4][10] ),
    .A1(_07211_),
    .S(_01654_),
    .X(_01655_));
 sky130_fd_sc_hd__buf_1 _14472_ (.A(_01655_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_2 _14473_ (.A0(\core.cpuregs[4][11] ),
    .A1(_07214_),
    .S(_01654_),
    .X(_01656_));
 sky130_fd_sc_hd__buf_1 _14474_ (.A(_01656_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_2 _14475_ (.A0(\core.cpuregs[4][12] ),
    .A1(_07216_),
    .S(_01654_),
    .X(_01657_));
 sky130_fd_sc_hd__buf_1 _14476_ (.A(_01657_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_2 _14477_ (.A0(\core.cpuregs[4][13] ),
    .A1(_07218_),
    .S(_01654_),
    .X(_01658_));
 sky130_fd_sc_hd__buf_1 _14478_ (.A(_01658_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_2 _14479_ (.A0(\core.cpuregs[4][14] ),
    .A1(_07220_),
    .S(_01654_),
    .X(_01659_));
 sky130_fd_sc_hd__buf_1 _14480_ (.A(_01659_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_2 _14481_ (.A0(\core.cpuregs[4][15] ),
    .A1(_07222_),
    .S(_01654_),
    .X(_01660_));
 sky130_fd_sc_hd__buf_1 _14482_ (.A(_01660_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_2 _14483_ (.A0(\core.cpuregs[4][16] ),
    .A1(_07224_),
    .S(_01654_),
    .X(_01661_));
 sky130_fd_sc_hd__buf_1 _14484_ (.A(_01661_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_2 _14485_ (.A0(\core.cpuregs[4][17] ),
    .A1(_07226_),
    .S(_01654_),
    .X(_01662_));
 sky130_fd_sc_hd__buf_1 _14486_ (.A(_01662_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_2 _14487_ (.A0(\core.cpuregs[4][18] ),
    .A1(_07228_),
    .S(_01654_),
    .X(_01663_));
 sky130_fd_sc_hd__buf_1 _14488_ (.A(_01663_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_2 _14489_ (.A0(\core.cpuregs[4][19] ),
    .A1(_07230_),
    .S(_01654_),
    .X(_01664_));
 sky130_fd_sc_hd__buf_1 _14490_ (.A(_01664_),
    .X(_01234_));
 sky130_fd_sc_hd__buf_1 _14491_ (.A(_01642_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_2 _14492_ (.A0(\core.cpuregs[4][20] ),
    .A1(_07232_),
    .S(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__buf_1 _14493_ (.A(_01666_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_2 _14494_ (.A0(\core.cpuregs[4][21] ),
    .A1(_07235_),
    .S(_01665_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_1 _14495_ (.A(_01667_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_2 _14496_ (.A0(\core.cpuregs[4][22] ),
    .A1(_07237_),
    .S(_01665_),
    .X(_01668_));
 sky130_fd_sc_hd__buf_1 _14497_ (.A(_01668_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_2 _14498_ (.A0(\core.cpuregs[4][23] ),
    .A1(_07239_),
    .S(_01665_),
    .X(_01669_));
 sky130_fd_sc_hd__buf_1 _14499_ (.A(_01669_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_2 _14500_ (.A0(\core.cpuregs[4][24] ),
    .A1(_07241_),
    .S(_01665_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_1 _14501_ (.A(_01670_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_2 _14502_ (.A0(\core.cpuregs[4][25] ),
    .A1(_07243_),
    .S(_01665_),
    .X(_01671_));
 sky130_fd_sc_hd__buf_1 _14503_ (.A(_01671_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_2 _14504_ (.A0(\core.cpuregs[4][26] ),
    .A1(_07245_),
    .S(_01665_),
    .X(_01672_));
 sky130_fd_sc_hd__buf_1 _14505_ (.A(_01672_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_2 _14506_ (.A0(\core.cpuregs[4][27] ),
    .A1(_07247_),
    .S(_01665_),
    .X(_01673_));
 sky130_fd_sc_hd__buf_1 _14507_ (.A(_01673_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_2 _14508_ (.A0(\core.cpuregs[4][28] ),
    .A1(_07249_),
    .S(_01665_),
    .X(_01674_));
 sky130_fd_sc_hd__buf_1 _14509_ (.A(_01674_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_2 _14510_ (.A0(\core.cpuregs[4][29] ),
    .A1(_07251_),
    .S(_01665_),
    .X(_01675_));
 sky130_fd_sc_hd__buf_1 _14511_ (.A(_01675_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_2 _14512_ (.A0(\core.cpuregs[4][30] ),
    .A1(_07253_),
    .S(_01642_),
    .X(_01676_));
 sky130_fd_sc_hd__buf_1 _14513_ (.A(_01676_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_2 _14514_ (.A0(\core.cpuregs[4][31] ),
    .A1(_07255_),
    .S(_01642_),
    .X(_01677_));
 sky130_fd_sc_hd__buf_1 _14515_ (.A(_01677_),
    .X(_01246_));
 sky130_fd_sc_hd__nor2_2 _14516_ (.A(_05286_),
    .B(_05620_),
    .Y(_01678_));
 sky130_fd_sc_hd__buf_1 _14517_ (.A(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_2 _14518_ (.A0(\core.cpuregs[3][0] ),
    .A1(_07188_),
    .S(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__buf_1 _14519_ (.A(_01680_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_2 _14520_ (.A0(\core.cpuregs[3][1] ),
    .A1(_07193_),
    .S(_01679_),
    .X(_01681_));
 sky130_fd_sc_hd__buf_1 _14521_ (.A(_01681_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_2 _14522_ (.A0(\core.cpuregs[3][2] ),
    .A1(_07195_),
    .S(_01679_),
    .X(_01682_));
 sky130_fd_sc_hd__buf_1 _14523_ (.A(_01682_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_2 _14524_ (.A0(\core.cpuregs[3][3] ),
    .A1(_07197_),
    .S(_01679_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_1 _14525_ (.A(_01683_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_2 _14526_ (.A0(\core.cpuregs[3][4] ),
    .A1(_07199_),
    .S(_01679_),
    .X(_01684_));
 sky130_fd_sc_hd__buf_1 _14527_ (.A(_01684_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_2 _14528_ (.A0(\core.cpuregs[3][5] ),
    .A1(_07201_),
    .S(_01679_),
    .X(_01685_));
 sky130_fd_sc_hd__buf_1 _14529_ (.A(_01685_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_2 _14530_ (.A0(\core.cpuregs[3][6] ),
    .A1(_07203_),
    .S(_01679_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_1 _14531_ (.A(_01686_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_2 _14532_ (.A0(\core.cpuregs[3][7] ),
    .A1(_07205_),
    .S(_01679_),
    .X(_01687_));
 sky130_fd_sc_hd__buf_1 _14533_ (.A(_01687_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_2 _14534_ (.A0(\core.cpuregs[3][8] ),
    .A1(_07207_),
    .S(_01679_),
    .X(_01688_));
 sky130_fd_sc_hd__buf_1 _14535_ (.A(_01688_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_2 _14536_ (.A0(\core.cpuregs[3][9] ),
    .A1(_07209_),
    .S(_01679_),
    .X(_01689_));
 sky130_fd_sc_hd__buf_1 _14537_ (.A(_01689_),
    .X(_01256_));
 sky130_fd_sc_hd__buf_1 _14538_ (.A(_01678_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_2 _14539_ (.A0(\core.cpuregs[3][10] ),
    .A1(_07211_),
    .S(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__buf_1 _14540_ (.A(_01691_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_2 _14541_ (.A0(\core.cpuregs[3][11] ),
    .A1(_07214_),
    .S(_01690_),
    .X(_01692_));
 sky130_fd_sc_hd__buf_1 _14542_ (.A(_01692_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_2 _14543_ (.A0(\core.cpuregs[3][12] ),
    .A1(_07216_),
    .S(_01690_),
    .X(_01693_));
 sky130_fd_sc_hd__buf_1 _14544_ (.A(_01693_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_2 _14545_ (.A0(\core.cpuregs[3][13] ),
    .A1(_07218_),
    .S(_01690_),
    .X(_01694_));
 sky130_fd_sc_hd__buf_1 _14546_ (.A(_01694_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_2 _14547_ (.A0(\core.cpuregs[3][14] ),
    .A1(_07220_),
    .S(_01690_),
    .X(_01695_));
 sky130_fd_sc_hd__buf_1 _14548_ (.A(_01695_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_2 _14549_ (.A0(\core.cpuregs[3][15] ),
    .A1(_07222_),
    .S(_01690_),
    .X(_01696_));
 sky130_fd_sc_hd__buf_1 _14550_ (.A(_01696_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_2 _14551_ (.A0(\core.cpuregs[3][16] ),
    .A1(_07224_),
    .S(_01690_),
    .X(_01697_));
 sky130_fd_sc_hd__buf_1 _14552_ (.A(_01697_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_2 _14553_ (.A0(\core.cpuregs[3][17] ),
    .A1(_07226_),
    .S(_01690_),
    .X(_01698_));
 sky130_fd_sc_hd__buf_1 _14554_ (.A(_01698_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_2 _14555_ (.A0(\core.cpuregs[3][18] ),
    .A1(_07228_),
    .S(_01690_),
    .X(_01699_));
 sky130_fd_sc_hd__buf_1 _14556_ (.A(_01699_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_2 _14557_ (.A0(\core.cpuregs[3][19] ),
    .A1(_07230_),
    .S(_01690_),
    .X(_01700_));
 sky130_fd_sc_hd__buf_1 _14558_ (.A(_01700_),
    .X(_01266_));
 sky130_fd_sc_hd__buf_1 _14559_ (.A(_01678_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_2 _14560_ (.A0(\core.cpuregs[3][20] ),
    .A1(_07232_),
    .S(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__buf_1 _14561_ (.A(_01702_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_2 _14562_ (.A0(\core.cpuregs[3][21] ),
    .A1(_07235_),
    .S(_01701_),
    .X(_01703_));
 sky130_fd_sc_hd__buf_1 _14563_ (.A(_01703_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_2 _14564_ (.A0(\core.cpuregs[3][22] ),
    .A1(_07237_),
    .S(_01701_),
    .X(_01704_));
 sky130_fd_sc_hd__buf_1 _14565_ (.A(_01704_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_2 _14566_ (.A0(\core.cpuregs[3][23] ),
    .A1(_07239_),
    .S(_01701_),
    .X(_01705_));
 sky130_fd_sc_hd__buf_1 _14567_ (.A(_01705_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_2 _14568_ (.A0(\core.cpuregs[3][24] ),
    .A1(_07241_),
    .S(_01701_),
    .X(_01706_));
 sky130_fd_sc_hd__buf_1 _14569_ (.A(_01706_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_2 _14570_ (.A0(\core.cpuregs[3][25] ),
    .A1(_07243_),
    .S(_01701_),
    .X(_01707_));
 sky130_fd_sc_hd__buf_1 _14571_ (.A(_01707_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_2 _14572_ (.A0(\core.cpuregs[3][26] ),
    .A1(_07245_),
    .S(_01701_),
    .X(_01708_));
 sky130_fd_sc_hd__buf_1 _14573_ (.A(_01708_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_2 _14574_ (.A0(\core.cpuregs[3][27] ),
    .A1(_07247_),
    .S(_01701_),
    .X(_01709_));
 sky130_fd_sc_hd__buf_1 _14575_ (.A(_01709_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_2 _14576_ (.A0(\core.cpuregs[3][28] ),
    .A1(_07249_),
    .S(_01701_),
    .X(_01710_));
 sky130_fd_sc_hd__buf_1 _14577_ (.A(_01710_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_2 _14578_ (.A0(\core.cpuregs[3][29] ),
    .A1(_07251_),
    .S(_01701_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_1 _14579_ (.A(_01711_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_2 _14580_ (.A0(\core.cpuregs[3][30] ),
    .A1(_07253_),
    .S(_01678_),
    .X(_01712_));
 sky130_fd_sc_hd__buf_1 _14581_ (.A(_01712_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_2 _14582_ (.A0(\core.cpuregs[3][31] ),
    .A1(_07255_),
    .S(_01678_),
    .X(_01713_));
 sky130_fd_sc_hd__buf_1 _14583_ (.A(_01713_),
    .X(_01278_));
 sky130_fd_sc_hd__nor2_2 _14584_ (.A(_05286_),
    .B(_07115_),
    .Y(_01714_));
 sky130_fd_sc_hd__buf_1 _14585_ (.A(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_2 _14586_ (.A0(\core.cpuregs[19][0] ),
    .A1(_07188_),
    .S(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__buf_1 _14587_ (.A(_01716_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_2 _14588_ (.A0(\core.cpuregs[19][1] ),
    .A1(_07193_),
    .S(_01715_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_1 _14589_ (.A(_01717_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_2 _14590_ (.A0(\core.cpuregs[19][2] ),
    .A1(_07195_),
    .S(_01715_),
    .X(_01718_));
 sky130_fd_sc_hd__buf_1 _14591_ (.A(_01718_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_2 _14592_ (.A0(\core.cpuregs[19][3] ),
    .A1(_07197_),
    .S(_01715_),
    .X(_01719_));
 sky130_fd_sc_hd__buf_1 _14593_ (.A(_01719_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_2 _14594_ (.A0(\core.cpuregs[19][4] ),
    .A1(_07199_),
    .S(_01715_),
    .X(_01720_));
 sky130_fd_sc_hd__buf_1 _14595_ (.A(_01720_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_2 _14596_ (.A0(\core.cpuregs[19][5] ),
    .A1(_07201_),
    .S(_01715_),
    .X(_01721_));
 sky130_fd_sc_hd__buf_1 _14597_ (.A(_01721_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_2 _14598_ (.A0(\core.cpuregs[19][6] ),
    .A1(_07203_),
    .S(_01715_),
    .X(_01722_));
 sky130_fd_sc_hd__buf_1 _14599_ (.A(_01722_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_2 _14600_ (.A0(\core.cpuregs[19][7] ),
    .A1(_07205_),
    .S(_01715_),
    .X(_01723_));
 sky130_fd_sc_hd__buf_1 _14601_ (.A(_01723_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_2 _14602_ (.A0(\core.cpuregs[19][8] ),
    .A1(_07207_),
    .S(_01715_),
    .X(_01724_));
 sky130_fd_sc_hd__buf_1 _14603_ (.A(_01724_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_2 _14604_ (.A0(\core.cpuregs[19][9] ),
    .A1(_07209_),
    .S(_01715_),
    .X(_01725_));
 sky130_fd_sc_hd__buf_1 _14605_ (.A(_01725_),
    .X(_01288_));
 sky130_fd_sc_hd__buf_1 _14606_ (.A(_01714_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_2 _14607_ (.A0(\core.cpuregs[19][10] ),
    .A1(_07211_),
    .S(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__buf_1 _14608_ (.A(_01727_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_2 _14609_ (.A0(\core.cpuregs[19][11] ),
    .A1(_07214_),
    .S(_01726_),
    .X(_01728_));
 sky130_fd_sc_hd__buf_1 _14610_ (.A(_01728_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_2 _14611_ (.A0(\core.cpuregs[19][12] ),
    .A1(_07216_),
    .S(_01726_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_1 _14612_ (.A(_01729_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_2 _14613_ (.A0(\core.cpuregs[19][13] ),
    .A1(_07218_),
    .S(_01726_),
    .X(_01730_));
 sky130_fd_sc_hd__buf_1 _14614_ (.A(_01730_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_2 _14615_ (.A0(\core.cpuregs[19][14] ),
    .A1(_07220_),
    .S(_01726_),
    .X(_01731_));
 sky130_fd_sc_hd__buf_1 _14616_ (.A(_01731_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_2 _14617_ (.A0(\core.cpuregs[19][15] ),
    .A1(_07222_),
    .S(_01726_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_1 _14618_ (.A(_01732_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_2 _14619_ (.A0(\core.cpuregs[19][16] ),
    .A1(_07224_),
    .S(_01726_),
    .X(_01733_));
 sky130_fd_sc_hd__buf_1 _14620_ (.A(_01733_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_2 _14621_ (.A0(\core.cpuregs[19][17] ),
    .A1(_07226_),
    .S(_01726_),
    .X(_01734_));
 sky130_fd_sc_hd__buf_1 _14622_ (.A(_01734_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_2 _14623_ (.A0(\core.cpuregs[19][18] ),
    .A1(_07228_),
    .S(_01726_),
    .X(_01735_));
 sky130_fd_sc_hd__buf_1 _14624_ (.A(_01735_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_2 _14625_ (.A0(\core.cpuregs[19][19] ),
    .A1(_07230_),
    .S(_01726_),
    .X(_01736_));
 sky130_fd_sc_hd__buf_1 _14626_ (.A(_01736_),
    .X(_01298_));
 sky130_fd_sc_hd__buf_1 _14627_ (.A(_01714_),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_2 _14628_ (.A0(\core.cpuregs[19][20] ),
    .A1(_07232_),
    .S(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__buf_1 _14629_ (.A(_01738_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_2 _14630_ (.A0(\core.cpuregs[19][21] ),
    .A1(_07235_),
    .S(_01737_),
    .X(_01739_));
 sky130_fd_sc_hd__buf_1 _14631_ (.A(_01739_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_2 _14632_ (.A0(\core.cpuregs[19][22] ),
    .A1(_07237_),
    .S(_01737_),
    .X(_01740_));
 sky130_fd_sc_hd__buf_1 _14633_ (.A(_01740_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_2 _14634_ (.A0(\core.cpuregs[19][23] ),
    .A1(_07239_),
    .S(_01737_),
    .X(_01741_));
 sky130_fd_sc_hd__buf_1 _14635_ (.A(_01741_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_2 _14636_ (.A0(\core.cpuregs[19][24] ),
    .A1(_07241_),
    .S(_01737_),
    .X(_01742_));
 sky130_fd_sc_hd__buf_1 _14637_ (.A(_01742_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_2 _14638_ (.A0(\core.cpuregs[19][25] ),
    .A1(_07243_),
    .S(_01737_),
    .X(_01743_));
 sky130_fd_sc_hd__buf_1 _14639_ (.A(_01743_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_2 _14640_ (.A0(\core.cpuregs[19][26] ),
    .A1(_07245_),
    .S(_01737_),
    .X(_01744_));
 sky130_fd_sc_hd__buf_1 _14641_ (.A(_01744_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_2 _14642_ (.A0(\core.cpuregs[19][27] ),
    .A1(_07247_),
    .S(_01737_),
    .X(_01745_));
 sky130_fd_sc_hd__buf_1 _14643_ (.A(_01745_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_2 _14644_ (.A0(\core.cpuregs[19][28] ),
    .A1(_07249_),
    .S(_01737_),
    .X(_01746_));
 sky130_fd_sc_hd__buf_1 _14645_ (.A(_01746_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_2 _14646_ (.A0(\core.cpuregs[19][29] ),
    .A1(_07251_),
    .S(_01737_),
    .X(_01747_));
 sky130_fd_sc_hd__buf_1 _14647_ (.A(_01747_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_2 _14648_ (.A0(\core.cpuregs[19][30] ),
    .A1(_07253_),
    .S(_01714_),
    .X(_01748_));
 sky130_fd_sc_hd__buf_1 _14649_ (.A(_01748_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_2 _14650_ (.A0(\core.cpuregs[19][31] ),
    .A1(_07255_),
    .S(_01714_),
    .X(_01749_));
 sky130_fd_sc_hd__buf_1 _14651_ (.A(_01749_),
    .X(_01310_));
 sky130_fd_sc_hd__nor2_2 _14652_ (.A(_05286_),
    .B(_05461_),
    .Y(_01750_));
 sky130_fd_sc_hd__buf_1 _14653_ (.A(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_2 _14654_ (.A0(\core.cpuregs[31][0] ),
    .A1(_07188_),
    .S(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__buf_1 _14655_ (.A(_01752_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_2 _14656_ (.A0(\core.cpuregs[31][1] ),
    .A1(_07193_),
    .S(_01751_),
    .X(_01753_));
 sky130_fd_sc_hd__buf_1 _14657_ (.A(_01753_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_2 _14658_ (.A0(\core.cpuregs[31][2] ),
    .A1(_07195_),
    .S(_01751_),
    .X(_01754_));
 sky130_fd_sc_hd__buf_1 _14659_ (.A(_01754_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_2 _14660_ (.A0(\core.cpuregs[31][3] ),
    .A1(_07197_),
    .S(_01751_),
    .X(_01755_));
 sky130_fd_sc_hd__buf_1 _14661_ (.A(_01755_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_2 _14662_ (.A0(\core.cpuregs[31][4] ),
    .A1(_07199_),
    .S(_01751_),
    .X(_01756_));
 sky130_fd_sc_hd__buf_1 _14663_ (.A(_01756_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_2 _14664_ (.A0(\core.cpuregs[31][5] ),
    .A1(_07201_),
    .S(_01751_),
    .X(_01757_));
 sky130_fd_sc_hd__buf_1 _14665_ (.A(_01757_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_2 _14666_ (.A0(\core.cpuregs[31][6] ),
    .A1(_07203_),
    .S(_01751_),
    .X(_01758_));
 sky130_fd_sc_hd__buf_1 _14667_ (.A(_01758_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_2 _14668_ (.A0(\core.cpuregs[31][7] ),
    .A1(_07205_),
    .S(_01751_),
    .X(_01759_));
 sky130_fd_sc_hd__buf_1 _14669_ (.A(_01759_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_2 _14670_ (.A0(\core.cpuregs[31][8] ),
    .A1(_07207_),
    .S(_01751_),
    .X(_01760_));
 sky130_fd_sc_hd__buf_1 _14671_ (.A(_01760_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_2 _14672_ (.A0(\core.cpuregs[31][9] ),
    .A1(_07209_),
    .S(_01751_),
    .X(_01761_));
 sky130_fd_sc_hd__buf_1 _14673_ (.A(_01761_),
    .X(_01320_));
 sky130_fd_sc_hd__buf_1 _14674_ (.A(_01750_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_2 _14675_ (.A0(\core.cpuregs[31][10] ),
    .A1(_07211_),
    .S(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__buf_1 _14676_ (.A(_01763_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_2 _14677_ (.A0(\core.cpuregs[31][11] ),
    .A1(_07214_),
    .S(_01762_),
    .X(_01764_));
 sky130_fd_sc_hd__buf_1 _14678_ (.A(_01764_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_2 _14679_ (.A0(\core.cpuregs[31][12] ),
    .A1(_07216_),
    .S(_01762_),
    .X(_01765_));
 sky130_fd_sc_hd__buf_1 _14680_ (.A(_01765_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_2 _14681_ (.A0(\core.cpuregs[31][13] ),
    .A1(_07218_),
    .S(_01762_),
    .X(_01766_));
 sky130_fd_sc_hd__buf_1 _14682_ (.A(_01766_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_2 _14683_ (.A0(\core.cpuregs[31][14] ),
    .A1(_07220_),
    .S(_01762_),
    .X(_01767_));
 sky130_fd_sc_hd__buf_1 _14684_ (.A(_01767_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_2 _14685_ (.A0(\core.cpuregs[31][15] ),
    .A1(_07222_),
    .S(_01762_),
    .X(_01768_));
 sky130_fd_sc_hd__buf_1 _14686_ (.A(_01768_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_2 _14687_ (.A0(\core.cpuregs[31][16] ),
    .A1(_07224_),
    .S(_01762_),
    .X(_01769_));
 sky130_fd_sc_hd__buf_1 _14688_ (.A(_01769_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_2 _14689_ (.A0(\core.cpuregs[31][17] ),
    .A1(_07226_),
    .S(_01762_),
    .X(_01770_));
 sky130_fd_sc_hd__buf_1 _14690_ (.A(_01770_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_2 _14691_ (.A0(\core.cpuregs[31][18] ),
    .A1(_07228_),
    .S(_01762_),
    .X(_01771_));
 sky130_fd_sc_hd__buf_1 _14692_ (.A(_01771_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_2 _14693_ (.A0(\core.cpuregs[31][19] ),
    .A1(_07230_),
    .S(_01762_),
    .X(_01772_));
 sky130_fd_sc_hd__buf_1 _14694_ (.A(_01772_),
    .X(_01330_));
 sky130_fd_sc_hd__buf_1 _14695_ (.A(_01750_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_2 _14696_ (.A0(\core.cpuregs[31][20] ),
    .A1(_07232_),
    .S(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__buf_1 _14697_ (.A(_01774_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_2 _14698_ (.A0(\core.cpuregs[31][21] ),
    .A1(_07235_),
    .S(_01773_),
    .X(_01775_));
 sky130_fd_sc_hd__buf_1 _14699_ (.A(_01775_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_2 _14700_ (.A0(\core.cpuregs[31][22] ),
    .A1(_07237_),
    .S(_01773_),
    .X(_01776_));
 sky130_fd_sc_hd__buf_1 _14701_ (.A(_01776_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_2 _14702_ (.A0(\core.cpuregs[31][23] ),
    .A1(_07239_),
    .S(_01773_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_1 _14703_ (.A(_01777_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_2 _14704_ (.A0(\core.cpuregs[31][24] ),
    .A1(_07241_),
    .S(_01773_),
    .X(_01778_));
 sky130_fd_sc_hd__buf_1 _14705_ (.A(_01778_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_2 _14706_ (.A0(\core.cpuregs[31][25] ),
    .A1(_07243_),
    .S(_01773_),
    .X(_01779_));
 sky130_fd_sc_hd__buf_1 _14707_ (.A(_01779_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_2 _14708_ (.A0(\core.cpuregs[31][26] ),
    .A1(_07245_),
    .S(_01773_),
    .X(_01780_));
 sky130_fd_sc_hd__buf_1 _14709_ (.A(_01780_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_2 _14710_ (.A0(\core.cpuregs[31][27] ),
    .A1(_07247_),
    .S(_01773_),
    .X(_01781_));
 sky130_fd_sc_hd__buf_1 _14711_ (.A(_01781_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_2 _14712_ (.A0(\core.cpuregs[31][28] ),
    .A1(_07249_),
    .S(_01773_),
    .X(_01782_));
 sky130_fd_sc_hd__buf_1 _14713_ (.A(_01782_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_2 _14714_ (.A0(\core.cpuregs[31][29] ),
    .A1(_07251_),
    .S(_01773_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_1 _14715_ (.A(_01783_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_2 _14716_ (.A0(\core.cpuregs[31][30] ),
    .A1(_07253_),
    .S(_01750_),
    .X(_01784_));
 sky130_fd_sc_hd__buf_1 _14717_ (.A(_01784_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_2 _14718_ (.A0(\core.cpuregs[31][31] ),
    .A1(_07255_),
    .S(_01750_),
    .X(_01785_));
 sky130_fd_sc_hd__buf_1 _14719_ (.A(_01785_),
    .X(_01342_));
 sky130_fd_sc_hd__nor2_2 _14720_ (.A(_05461_),
    .B(_05837_),
    .Y(_01786_));
 sky130_fd_sc_hd__buf_1 _14721_ (.A(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_2 _14722_ (.A0(\core.cpuregs[29][0] ),
    .A1(_07188_),
    .S(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__buf_1 _14723_ (.A(_01788_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_2 _14724_ (.A0(\core.cpuregs[29][1] ),
    .A1(_07193_),
    .S(_01787_),
    .X(_01789_));
 sky130_fd_sc_hd__buf_1 _14725_ (.A(_01789_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_2 _14726_ (.A0(\core.cpuregs[29][2] ),
    .A1(_07195_),
    .S(_01787_),
    .X(_01790_));
 sky130_fd_sc_hd__buf_1 _14727_ (.A(_01790_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_2 _14728_ (.A0(\core.cpuregs[29][3] ),
    .A1(_07197_),
    .S(_01787_),
    .X(_01791_));
 sky130_fd_sc_hd__buf_1 _14729_ (.A(_01791_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_2 _14730_ (.A0(\core.cpuregs[29][4] ),
    .A1(_07199_),
    .S(_01787_),
    .X(_01792_));
 sky130_fd_sc_hd__buf_1 _14731_ (.A(_01792_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_2 _14732_ (.A0(\core.cpuregs[29][5] ),
    .A1(_07201_),
    .S(_01787_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_1 _14733_ (.A(_01793_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_2 _14734_ (.A0(\core.cpuregs[29][6] ),
    .A1(_07203_),
    .S(_01787_),
    .X(_01794_));
 sky130_fd_sc_hd__buf_1 _14735_ (.A(_01794_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_2 _14736_ (.A0(\core.cpuregs[29][7] ),
    .A1(_07205_),
    .S(_01787_),
    .X(_01795_));
 sky130_fd_sc_hd__buf_1 _14737_ (.A(_01795_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_2 _14738_ (.A0(\core.cpuregs[29][8] ),
    .A1(_07207_),
    .S(_01787_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_1 _14739_ (.A(_01796_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_2 _14740_ (.A0(\core.cpuregs[29][9] ),
    .A1(_07209_),
    .S(_01787_),
    .X(_01797_));
 sky130_fd_sc_hd__buf_1 _14741_ (.A(_01797_),
    .X(_01384_));
 sky130_fd_sc_hd__buf_1 _14742_ (.A(_01786_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_2 _14743_ (.A0(\core.cpuregs[29][10] ),
    .A1(_07211_),
    .S(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__buf_1 _14744_ (.A(_01799_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_2 _14745_ (.A0(\core.cpuregs[29][11] ),
    .A1(_07214_),
    .S(_01798_),
    .X(_01800_));
 sky130_fd_sc_hd__buf_1 _14746_ (.A(_01800_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_2 _14747_ (.A0(\core.cpuregs[29][12] ),
    .A1(_07216_),
    .S(_01798_),
    .X(_01801_));
 sky130_fd_sc_hd__buf_1 _14748_ (.A(_01801_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_2 _14749_ (.A0(\core.cpuregs[29][13] ),
    .A1(_07218_),
    .S(_01798_),
    .X(_01802_));
 sky130_fd_sc_hd__buf_1 _14750_ (.A(_01802_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_2 _14751_ (.A0(\core.cpuregs[29][14] ),
    .A1(_07220_),
    .S(_01798_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _14752_ (.A(_01803_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_2 _14753_ (.A0(\core.cpuregs[29][15] ),
    .A1(_07222_),
    .S(_01798_),
    .X(_01804_));
 sky130_fd_sc_hd__buf_1 _14754_ (.A(_01804_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_2 _14755_ (.A0(\core.cpuregs[29][16] ),
    .A1(_07224_),
    .S(_01798_),
    .X(_01805_));
 sky130_fd_sc_hd__buf_1 _14756_ (.A(_01805_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_2 _14757_ (.A0(\core.cpuregs[29][17] ),
    .A1(_07226_),
    .S(_01798_),
    .X(_01806_));
 sky130_fd_sc_hd__buf_1 _14758_ (.A(_01806_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_2 _14759_ (.A0(\core.cpuregs[29][18] ),
    .A1(_07228_),
    .S(_01798_),
    .X(_01807_));
 sky130_fd_sc_hd__buf_1 _14760_ (.A(_01807_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_2 _14761_ (.A0(\core.cpuregs[29][19] ),
    .A1(_07230_),
    .S(_01798_),
    .X(_01808_));
 sky130_fd_sc_hd__buf_1 _14762_ (.A(_01808_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_1 _14763_ (.A(_01786_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_2 _14764_ (.A0(\core.cpuregs[29][20] ),
    .A1(_07232_),
    .S(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__buf_1 _14765_ (.A(_01810_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_2 _14766_ (.A0(\core.cpuregs[29][21] ),
    .A1(_07235_),
    .S(_01809_),
    .X(_01811_));
 sky130_fd_sc_hd__buf_1 _14767_ (.A(_01811_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_2 _14768_ (.A0(\core.cpuregs[29][22] ),
    .A1(_07237_),
    .S(_01809_),
    .X(_01812_));
 sky130_fd_sc_hd__buf_1 _14769_ (.A(_01812_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_2 _14770_ (.A0(\core.cpuregs[29][23] ),
    .A1(_07239_),
    .S(_01809_),
    .X(_01813_));
 sky130_fd_sc_hd__buf_1 _14771_ (.A(_01813_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_2 _14772_ (.A0(\core.cpuregs[29][24] ),
    .A1(_07241_),
    .S(_01809_),
    .X(_01814_));
 sky130_fd_sc_hd__buf_1 _14773_ (.A(_01814_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_2 _14774_ (.A0(\core.cpuregs[29][25] ),
    .A1(_07243_),
    .S(_01809_),
    .X(_01815_));
 sky130_fd_sc_hd__buf_1 _14775_ (.A(_01815_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_2 _14776_ (.A0(\core.cpuregs[29][26] ),
    .A1(_07245_),
    .S(_01809_),
    .X(_01816_));
 sky130_fd_sc_hd__buf_1 _14777_ (.A(_01816_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_2 _14778_ (.A0(\core.cpuregs[29][27] ),
    .A1(_07247_),
    .S(_01809_),
    .X(_01817_));
 sky130_fd_sc_hd__buf_1 _14779_ (.A(_01817_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_2 _14780_ (.A0(\core.cpuregs[29][28] ),
    .A1(_07249_),
    .S(_01809_),
    .X(_01818_));
 sky130_fd_sc_hd__buf_1 _14781_ (.A(_01818_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_2 _14782_ (.A0(\core.cpuregs[29][29] ),
    .A1(_07251_),
    .S(_01809_),
    .X(_01819_));
 sky130_fd_sc_hd__buf_1 _14783_ (.A(_01819_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_2 _14784_ (.A0(\core.cpuregs[29][30] ),
    .A1(_07253_),
    .S(_01786_),
    .X(_01820_));
 sky130_fd_sc_hd__buf_1 _14785_ (.A(_01820_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_2 _14786_ (.A0(\core.cpuregs[29][31] ),
    .A1(_07255_),
    .S(_01786_),
    .X(_01821_));
 sky130_fd_sc_hd__buf_1 _14787_ (.A(_01821_),
    .X(_01406_));
 sky130_fd_sc_hd__or2_2 _14788_ (.A(_05464_),
    .B(_07115_),
    .X(_01822_));
 sky130_fd_sc_hd__buf_1 _14789_ (.A(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_2 _14790_ (.A0(_05284_),
    .A1(\core.cpuregs[18][0] ),
    .S(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__buf_1 _14791_ (.A(_01824_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_2 _14792_ (.A0(_05292_),
    .A1(\core.cpuregs[18][1] ),
    .S(_01823_),
    .X(_01825_));
 sky130_fd_sc_hd__buf_1 _14793_ (.A(_01825_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_2 _14794_ (.A0(_05297_),
    .A1(\core.cpuregs[18][2] ),
    .S(_01823_),
    .X(_01826_));
 sky130_fd_sc_hd__buf_1 _14795_ (.A(_01826_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_2 _14796_ (.A0(_05304_),
    .A1(\core.cpuregs[18][3] ),
    .S(_01823_),
    .X(_01827_));
 sky130_fd_sc_hd__buf_1 _14797_ (.A(_01827_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_2 _14798_ (.A0(_05310_),
    .A1(\core.cpuregs[18][4] ),
    .S(_01823_),
    .X(_01828_));
 sky130_fd_sc_hd__buf_1 _14799_ (.A(_01828_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_2 _14800_ (.A0(_05315_),
    .A1(\core.cpuregs[18][5] ),
    .S(_01823_),
    .X(_01829_));
 sky130_fd_sc_hd__buf_1 _14801_ (.A(_01829_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_2 _14802_ (.A0(_05320_),
    .A1(\core.cpuregs[18][6] ),
    .S(_01823_),
    .X(_01830_));
 sky130_fd_sc_hd__buf_1 _14803_ (.A(_01830_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_2 _14804_ (.A0(_05326_),
    .A1(\core.cpuregs[18][7] ),
    .S(_01823_),
    .X(_01831_));
 sky130_fd_sc_hd__buf_1 _14805_ (.A(_01831_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_2 _14806_ (.A0(_05332_),
    .A1(\core.cpuregs[18][8] ),
    .S(_01823_),
    .X(_01832_));
 sky130_fd_sc_hd__buf_1 _14807_ (.A(_01832_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_2 _14808_ (.A0(_05337_),
    .A1(\core.cpuregs[18][9] ),
    .S(_01823_),
    .X(_01833_));
 sky130_fd_sc_hd__buf_1 _14809_ (.A(_01833_),
    .X(_01416_));
 sky130_fd_sc_hd__buf_1 _14810_ (.A(_01822_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_2 _14811_ (.A0(_05343_),
    .A1(\core.cpuregs[18][10] ),
    .S(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__buf_1 _14812_ (.A(_01835_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_2 _14813_ (.A0(_05349_),
    .A1(\core.cpuregs[18][11] ),
    .S(_01834_),
    .X(_01836_));
 sky130_fd_sc_hd__buf_1 _14814_ (.A(_01836_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_2 _14815_ (.A0(_05355_),
    .A1(\core.cpuregs[18][12] ),
    .S(_01834_),
    .X(_01837_));
 sky130_fd_sc_hd__buf_1 _14816_ (.A(_01837_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_2 _14817_ (.A0(_05360_),
    .A1(\core.cpuregs[18][13] ),
    .S(_01834_),
    .X(_01838_));
 sky130_fd_sc_hd__buf_1 _14818_ (.A(_01838_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_2 _14819_ (.A0(_05367_),
    .A1(\core.cpuregs[18][14] ),
    .S(_01834_),
    .X(_01839_));
 sky130_fd_sc_hd__buf_1 _14820_ (.A(_01839_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_2 _14821_ (.A0(_05372_),
    .A1(\core.cpuregs[18][15] ),
    .S(_01834_),
    .X(_01840_));
 sky130_fd_sc_hd__buf_1 _14822_ (.A(_01840_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_2 _14823_ (.A0(_05377_),
    .A1(\core.cpuregs[18][16] ),
    .S(_01834_),
    .X(_01841_));
 sky130_fd_sc_hd__buf_1 _14824_ (.A(_01841_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_2 _14825_ (.A0(_05383_),
    .A1(\core.cpuregs[18][17] ),
    .S(_01834_),
    .X(_01842_));
 sky130_fd_sc_hd__buf_1 _14826_ (.A(_01842_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_2 _14827_ (.A0(_05388_),
    .A1(\core.cpuregs[18][18] ),
    .S(_01834_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_1 _14828_ (.A(_01843_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_2 _14829_ (.A0(_05393_),
    .A1(\core.cpuregs[18][19] ),
    .S(_01834_),
    .X(_01844_));
 sky130_fd_sc_hd__buf_1 _14830_ (.A(_01844_),
    .X(_01426_));
 sky130_fd_sc_hd__buf_1 _14831_ (.A(_01822_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_2 _14832_ (.A0(_05399_),
    .A1(\core.cpuregs[18][20] ),
    .S(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__buf_1 _14833_ (.A(_01846_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_2 _14834_ (.A0(_05405_),
    .A1(\core.cpuregs[18][21] ),
    .S(_01845_),
    .X(_01847_));
 sky130_fd_sc_hd__buf_1 _14835_ (.A(_01847_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_2 _14836_ (.A0(_05410_),
    .A1(\core.cpuregs[18][22] ),
    .S(_01845_),
    .X(_01848_));
 sky130_fd_sc_hd__buf_1 _14837_ (.A(_01848_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_2 _14838_ (.A0(_05416_),
    .A1(\core.cpuregs[18][23] ),
    .S(_01845_),
    .X(_01849_));
 sky130_fd_sc_hd__buf_1 _14839_ (.A(_01849_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_2 _14840_ (.A0(_05421_),
    .A1(\core.cpuregs[18][24] ),
    .S(_01845_),
    .X(_01850_));
 sky130_fd_sc_hd__buf_1 _14841_ (.A(_01850_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_2 _14842_ (.A0(_05426_),
    .A1(\core.cpuregs[18][25] ),
    .S(_01845_),
    .X(_01851_));
 sky130_fd_sc_hd__buf_1 _14843_ (.A(_01851_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_2 _14844_ (.A0(_05432_),
    .A1(\core.cpuregs[18][26] ),
    .S(_01845_),
    .X(_01852_));
 sky130_fd_sc_hd__buf_1 _14845_ (.A(_01852_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_2 _14846_ (.A0(_05437_),
    .A1(\core.cpuregs[18][27] ),
    .S(_01845_),
    .X(_01853_));
 sky130_fd_sc_hd__buf_1 _14847_ (.A(_01853_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_2 _14848_ (.A0(_05442_),
    .A1(\core.cpuregs[18][28] ),
    .S(_01845_),
    .X(_01854_));
 sky130_fd_sc_hd__buf_1 _14849_ (.A(_01854_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_2 _14850_ (.A0(_05448_),
    .A1(\core.cpuregs[18][29] ),
    .S(_01845_),
    .X(_01855_));
 sky130_fd_sc_hd__buf_1 _14851_ (.A(_01855_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_2 _14852_ (.A0(_05453_),
    .A1(\core.cpuregs[18][30] ),
    .S(_01822_),
    .X(_01856_));
 sky130_fd_sc_hd__buf_1 _14853_ (.A(_01856_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_2 _14854_ (.A0(_05458_),
    .A1(\core.cpuregs[18][31] ),
    .S(_01822_),
    .X(_01857_));
 sky130_fd_sc_hd__buf_1 _14855_ (.A(_01857_),
    .X(_01438_));
 sky130_fd_sc_hd__nor2_2 _14856_ (.A(_05657_),
    .B(_05766_),
    .Y(_01858_));
 sky130_fd_sc_hd__buf_1 _14857_ (.A(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_2 _14858_ (.A0(\core.cpuregs[24][0] ),
    .A1(_05283_),
    .S(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_1 _14859_ (.A(_01860_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_2 _14860_ (.A0(\core.cpuregs[24][1] ),
    .A1(_05291_),
    .S(_01859_),
    .X(_01861_));
 sky130_fd_sc_hd__buf_1 _14861_ (.A(_01861_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_2 _14862_ (.A0(\core.cpuregs[24][2] ),
    .A1(_05296_),
    .S(_01859_),
    .X(_01862_));
 sky130_fd_sc_hd__buf_1 _14863_ (.A(_01862_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_2 _14864_ (.A0(\core.cpuregs[24][3] ),
    .A1(_05303_),
    .S(_01859_),
    .X(_01863_));
 sky130_fd_sc_hd__buf_1 _14865_ (.A(_01863_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_2 _14866_ (.A0(\core.cpuregs[24][4] ),
    .A1(_05309_),
    .S(_01859_),
    .X(_01864_));
 sky130_fd_sc_hd__buf_1 _14867_ (.A(_01864_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_2 _14868_ (.A0(\core.cpuregs[24][5] ),
    .A1(_05314_),
    .S(_01859_),
    .X(_01865_));
 sky130_fd_sc_hd__buf_1 _14869_ (.A(_01865_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_2 _14870_ (.A0(\core.cpuregs[24][6] ),
    .A1(_05319_),
    .S(_01859_),
    .X(_01866_));
 sky130_fd_sc_hd__buf_1 _14871_ (.A(_01866_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_2 _14872_ (.A0(\core.cpuregs[24][7] ),
    .A1(_05325_),
    .S(_01859_),
    .X(_01867_));
 sky130_fd_sc_hd__buf_1 _14873_ (.A(_01867_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_2 _14874_ (.A0(\core.cpuregs[24][8] ),
    .A1(_05331_),
    .S(_01859_),
    .X(_01868_));
 sky130_fd_sc_hd__buf_1 _14875_ (.A(_01868_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_2 _14876_ (.A0(\core.cpuregs[24][9] ),
    .A1(_05336_),
    .S(_01859_),
    .X(_01869_));
 sky130_fd_sc_hd__buf_1 _14877_ (.A(_01869_),
    .X(_01448_));
 sky130_fd_sc_hd__buf_1 _14878_ (.A(_01858_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_2 _14879_ (.A0(\core.cpuregs[24][10] ),
    .A1(_05342_),
    .S(_01870_),
    .X(_01871_));
 sky130_fd_sc_hd__buf_1 _14880_ (.A(_01871_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_2 _14881_ (.A0(\core.cpuregs[24][11] ),
    .A1(_05348_),
    .S(_01870_),
    .X(_01872_));
 sky130_fd_sc_hd__buf_1 _14882_ (.A(_01872_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_2 _14883_ (.A0(\core.cpuregs[24][12] ),
    .A1(_05354_),
    .S(_01870_),
    .X(_01873_));
 sky130_fd_sc_hd__buf_1 _14884_ (.A(_01873_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_2 _14885_ (.A0(\core.cpuregs[24][13] ),
    .A1(_05359_),
    .S(_01870_),
    .X(_01874_));
 sky130_fd_sc_hd__buf_1 _14886_ (.A(_01874_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_2 _14887_ (.A0(\core.cpuregs[24][14] ),
    .A1(_05366_),
    .S(_01870_),
    .X(_01875_));
 sky130_fd_sc_hd__buf_1 _14888_ (.A(_01875_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_2 _14889_ (.A0(\core.cpuregs[24][15] ),
    .A1(_05371_),
    .S(_01870_),
    .X(_01876_));
 sky130_fd_sc_hd__buf_1 _14890_ (.A(_01876_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_2 _14891_ (.A0(\core.cpuregs[24][16] ),
    .A1(_05376_),
    .S(_01870_),
    .X(_01877_));
 sky130_fd_sc_hd__buf_1 _14892_ (.A(_01877_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_2 _14893_ (.A0(\core.cpuregs[24][17] ),
    .A1(_05382_),
    .S(_01870_),
    .X(_01878_));
 sky130_fd_sc_hd__buf_1 _14894_ (.A(_01878_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_2 _14895_ (.A0(\core.cpuregs[24][18] ),
    .A1(_05387_),
    .S(_01870_),
    .X(_01879_));
 sky130_fd_sc_hd__buf_1 _14896_ (.A(_01879_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_2 _14897_ (.A0(\core.cpuregs[24][19] ),
    .A1(_05392_),
    .S(_01870_),
    .X(_01880_));
 sky130_fd_sc_hd__buf_1 _14898_ (.A(_01880_),
    .X(_01458_));
 sky130_fd_sc_hd__buf_1 _14899_ (.A(_01858_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_2 _14900_ (.A0(\core.cpuregs[24][20] ),
    .A1(_05398_),
    .S(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_1 _14901_ (.A(_01882_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_2 _14902_ (.A0(\core.cpuregs[24][21] ),
    .A1(_05404_),
    .S(_01881_),
    .X(_01883_));
 sky130_fd_sc_hd__buf_1 _14903_ (.A(_01883_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_2 _14904_ (.A0(\core.cpuregs[24][22] ),
    .A1(_05409_),
    .S(_01881_),
    .X(_01884_));
 sky130_fd_sc_hd__buf_1 _14905_ (.A(_01884_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_2 _14906_ (.A0(\core.cpuregs[24][23] ),
    .A1(_05415_),
    .S(_01881_),
    .X(_01885_));
 sky130_fd_sc_hd__buf_1 _14907_ (.A(_01885_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_2 _14908_ (.A0(\core.cpuregs[24][24] ),
    .A1(_05420_),
    .S(_01881_),
    .X(_01886_));
 sky130_fd_sc_hd__buf_1 _14909_ (.A(_01886_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_2 _14910_ (.A0(\core.cpuregs[24][25] ),
    .A1(_05425_),
    .S(_01881_),
    .X(_01887_));
 sky130_fd_sc_hd__buf_1 _14911_ (.A(_01887_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_2 _14912_ (.A0(\core.cpuregs[24][26] ),
    .A1(_05431_),
    .S(_01881_),
    .X(_01888_));
 sky130_fd_sc_hd__buf_1 _14913_ (.A(_01888_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_2 _14914_ (.A0(\core.cpuregs[24][27] ),
    .A1(_05436_),
    .S(_01881_),
    .X(_01889_));
 sky130_fd_sc_hd__buf_1 _14915_ (.A(_01889_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_2 _14916_ (.A0(\core.cpuregs[24][28] ),
    .A1(_05441_),
    .S(_01881_),
    .X(_01890_));
 sky130_fd_sc_hd__buf_1 _14917_ (.A(_01890_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_2 _14918_ (.A0(\core.cpuregs[24][29] ),
    .A1(_05447_),
    .S(_01881_),
    .X(_01891_));
 sky130_fd_sc_hd__buf_1 _14919_ (.A(_01891_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_2 _14920_ (.A0(\core.cpuregs[24][30] ),
    .A1(_05452_),
    .S(_01858_),
    .X(_01892_));
 sky130_fd_sc_hd__buf_1 _14921_ (.A(_01892_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_2 _14922_ (.A0(\core.cpuregs[24][31] ),
    .A1(_05457_),
    .S(_01858_),
    .X(_01893_));
 sky130_fd_sc_hd__buf_1 _14923_ (.A(_01893_),
    .X(_01470_));
 sky130_fd_sc_hd__or2_2 _14924_ (.A(_05837_),
    .B(_07365_),
    .X(_01894_));
 sky130_fd_sc_hd__buf_1 _14925_ (.A(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_2 _14926_ (.A0(_05284_),
    .A1(\core.cpuregs[9][0] ),
    .S(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__buf_1 _14927_ (.A(_01896_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_2 _14928_ (.A0(_05292_),
    .A1(\core.cpuregs[9][1] ),
    .S(_01895_),
    .X(_01897_));
 sky130_fd_sc_hd__buf_1 _14929_ (.A(_01897_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_2 _14930_ (.A0(_05297_),
    .A1(\core.cpuregs[9][2] ),
    .S(_01895_),
    .X(_01898_));
 sky130_fd_sc_hd__buf_1 _14931_ (.A(_01898_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_2 _14932_ (.A0(_05304_),
    .A1(\core.cpuregs[9][3] ),
    .S(_01895_),
    .X(_01899_));
 sky130_fd_sc_hd__buf_1 _14933_ (.A(_01899_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_2 _14934_ (.A0(_05310_),
    .A1(\core.cpuregs[9][4] ),
    .S(_01895_),
    .X(_01900_));
 sky130_fd_sc_hd__buf_1 _14935_ (.A(_01900_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_2 _14936_ (.A0(_05315_),
    .A1(\core.cpuregs[9][5] ),
    .S(_01895_),
    .X(_01901_));
 sky130_fd_sc_hd__buf_1 _14937_ (.A(_01901_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_2 _14938_ (.A0(_05320_),
    .A1(\core.cpuregs[9][6] ),
    .S(_01895_),
    .X(_01902_));
 sky130_fd_sc_hd__buf_1 _14939_ (.A(_01902_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_2 _14940_ (.A0(_05326_),
    .A1(\core.cpuregs[9][7] ),
    .S(_01895_),
    .X(_01903_));
 sky130_fd_sc_hd__buf_1 _14941_ (.A(_01903_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_2 _14942_ (.A0(_05332_),
    .A1(\core.cpuregs[9][8] ),
    .S(_01895_),
    .X(_01904_));
 sky130_fd_sc_hd__buf_1 _14943_ (.A(_01904_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_2 _14944_ (.A0(_05337_),
    .A1(\core.cpuregs[9][9] ),
    .S(_01895_),
    .X(_01905_));
 sky130_fd_sc_hd__buf_1 _14945_ (.A(_01905_),
    .X(_01480_));
 sky130_fd_sc_hd__buf_1 _14946_ (.A(_01894_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_2 _14947_ (.A0(_05343_),
    .A1(\core.cpuregs[9][10] ),
    .S(_01906_),
    .X(_01907_));
 sky130_fd_sc_hd__buf_1 _14948_ (.A(_01907_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_2 _14949_ (.A0(_05349_),
    .A1(\core.cpuregs[9][11] ),
    .S(_01906_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_1 _14950_ (.A(_01908_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_2 _14951_ (.A0(_05355_),
    .A1(\core.cpuregs[9][12] ),
    .S(_01906_),
    .X(_01909_));
 sky130_fd_sc_hd__buf_1 _14952_ (.A(_01909_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_2 _14953_ (.A0(_05360_),
    .A1(\core.cpuregs[9][13] ),
    .S(_01906_),
    .X(_01910_));
 sky130_fd_sc_hd__buf_1 _14954_ (.A(_01910_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_2 _14955_ (.A0(_05367_),
    .A1(\core.cpuregs[9][14] ),
    .S(_01906_),
    .X(_01911_));
 sky130_fd_sc_hd__buf_1 _14956_ (.A(_01911_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_2 _14957_ (.A0(_05372_),
    .A1(\core.cpuregs[9][15] ),
    .S(_01906_),
    .X(_01912_));
 sky130_fd_sc_hd__buf_1 _14958_ (.A(_01912_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_2 _14959_ (.A0(_05377_),
    .A1(\core.cpuregs[9][16] ),
    .S(_01906_),
    .X(_01913_));
 sky130_fd_sc_hd__buf_1 _14960_ (.A(_01913_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_2 _14961_ (.A0(_05383_),
    .A1(\core.cpuregs[9][17] ),
    .S(_01906_),
    .X(_01914_));
 sky130_fd_sc_hd__buf_1 _14962_ (.A(_01914_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_2 _14963_ (.A0(_05388_),
    .A1(\core.cpuregs[9][18] ),
    .S(_01906_),
    .X(_01915_));
 sky130_fd_sc_hd__buf_1 _14964_ (.A(_01915_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_2 _14965_ (.A0(_05393_),
    .A1(\core.cpuregs[9][19] ),
    .S(_01906_),
    .X(_01916_));
 sky130_fd_sc_hd__buf_1 _14966_ (.A(_01916_),
    .X(_01490_));
 sky130_fd_sc_hd__buf_1 _14967_ (.A(_01894_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_2 _14968_ (.A0(_05399_),
    .A1(\core.cpuregs[9][20] ),
    .S(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__buf_1 _14969_ (.A(_01918_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_2 _14970_ (.A0(_05405_),
    .A1(\core.cpuregs[9][21] ),
    .S(_01917_),
    .X(_01919_));
 sky130_fd_sc_hd__buf_1 _14971_ (.A(_01919_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_2 _14972_ (.A0(_05410_),
    .A1(\core.cpuregs[9][22] ),
    .S(_01917_),
    .X(_01920_));
 sky130_fd_sc_hd__buf_1 _14973_ (.A(_01920_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_2 _14974_ (.A0(_05416_),
    .A1(\core.cpuregs[9][23] ),
    .S(_01917_),
    .X(_01921_));
 sky130_fd_sc_hd__buf_1 _14975_ (.A(_01921_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_2 _14976_ (.A0(_05421_),
    .A1(\core.cpuregs[9][24] ),
    .S(_01917_),
    .X(_01922_));
 sky130_fd_sc_hd__buf_1 _14977_ (.A(_01922_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_2 _14978_ (.A0(_05426_),
    .A1(\core.cpuregs[9][25] ),
    .S(_01917_),
    .X(_01923_));
 sky130_fd_sc_hd__buf_1 _14979_ (.A(_01923_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_2 _14980_ (.A0(_05432_),
    .A1(\core.cpuregs[9][26] ),
    .S(_01917_),
    .X(_01924_));
 sky130_fd_sc_hd__buf_1 _14981_ (.A(_01924_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_2 _14982_ (.A0(_05437_),
    .A1(\core.cpuregs[9][27] ),
    .S(_01917_),
    .X(_01925_));
 sky130_fd_sc_hd__buf_1 _14983_ (.A(_01925_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_2 _14984_ (.A0(_05442_),
    .A1(\core.cpuregs[9][28] ),
    .S(_01917_),
    .X(_01926_));
 sky130_fd_sc_hd__buf_1 _14985_ (.A(_01926_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_2 _14986_ (.A0(_05448_),
    .A1(\core.cpuregs[9][29] ),
    .S(_01917_),
    .X(_01927_));
 sky130_fd_sc_hd__buf_1 _14987_ (.A(_01927_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_2 _14988_ (.A0(_05453_),
    .A1(\core.cpuregs[9][30] ),
    .S(_01894_),
    .X(_01928_));
 sky130_fd_sc_hd__buf_1 _14989_ (.A(_01928_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_2 _14990_ (.A0(_05458_),
    .A1(\core.cpuregs[9][31] ),
    .S(_01894_),
    .X(_01929_));
 sky130_fd_sc_hd__buf_1 _14991_ (.A(_01929_),
    .X(_01502_));
 sky130_fd_sc_hd__a22o_2 _14992_ (.A1(\core.instr_lhu ),
    .A2(_05921_),
    .B1(_06900_),
    .B2(_02091_),
    .X(_01503_));
 sky130_fd_sc_hd__nor2_2 _14993_ (.A(_05830_),
    .B(_05950_),
    .Y(_01930_));
 sky130_fd_sc_hd__a22o_2 _14994_ (.A1(\core.instr_lbu ),
    .A2(_05921_),
    .B1(_01930_),
    .B2(_02091_),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_2 _14995_ (.A(_05943_),
    .B(_05922_),
    .Y(_01931_));
 sky130_fd_sc_hd__a22o_2 _14996_ (.A1(\core.instr_lw ),
    .A2(_05921_),
    .B1(_01931_),
    .B2(_02091_),
    .X(_01505_));
 sky130_fd_sc_hd__a22o_2 _14997_ (.A1(\core.instr_lh ),
    .A2(_05921_),
    .B1(_05833_),
    .B2(_02091_),
    .X(_01506_));
 sky130_fd_sc_hd__and3_2 _14998_ (.A(\core.mem_rdata_q[12] ),
    .B(\core.mem_rdata_q[13] ),
    .C(\core.mem_rdata_q[14] ),
    .X(_01932_));
 sky130_fd_sc_hd__a22o_2 _14999_ (.A1(\core.instr_bgeu ),
    .A2(_05932_),
    .B1(_06903_),
    .B2(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__and2_2 _15000_ (.A(_05928_),
    .B(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__buf_1 _15001_ (.A(_01934_),
    .X(_01507_));
 sky130_fd_sc_hd__a22o_2 _15002_ (.A1(\core.instr_blt ),
    .A2(_05932_),
    .B1(_01930_),
    .B2(\core.is_beq_bne_blt_bge_bltu_bgeu ),
    .X(_01935_));
 sky130_fd_sc_hd__and2_2 _15003_ (.A(_05928_),
    .B(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__buf_1 _15004_ (.A(_01936_),
    .X(_01508_));
 sky130_fd_sc_hd__and4bb_2 _15005_ (.A_N(\core.mem_rdata_q[20] ),
    .B_N(_05970_),
    .C(_05977_),
    .D(\core.mem_rdata_q[21] ),
    .X(_01937_));
 sky130_fd_sc_hd__a22o_2 _15006_ (.A1(_02456_),
    .A2(_05921_),
    .B1(_05969_),
    .B2(_01937_),
    .X(_01509_));
 sky130_fd_sc_hd__nor2_2 _15007_ (.A(\core.mem_rdata_q[24] ),
    .B(_05939_),
    .Y(_01938_));
 sky130_fd_sc_hd__a22o_2 _15008_ (.A1(_02684_),
    .A2(_05943_),
    .B1(_01937_),
    .B2(_01938_),
    .X(_01510_));
 sky130_fd_sc_hd__a32o_2 _15009_ (.A1(_05971_),
    .A2(_05977_),
    .A3(_01938_),
    .B1(_05943_),
    .B2(\core.instr_rdcycle ),
    .X(_01511_));
 sky130_fd_sc_hd__a22o_2 _15010_ (.A1(\core.instr_srai ),
    .A2(_05943_),
    .B1(_05925_),
    .B2(_05954_),
    .X(_01512_));
 sky130_fd_sc_hd__a22o_2 _15011_ (.A1(\core.instr_and ),
    .A2(_05932_),
    .B1(_05945_),
    .B2(_01932_),
    .X(_01939_));
 sky130_fd_sc_hd__and2_2 _15012_ (.A(_03546_),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__buf_1 _15013_ (.A(_01940_),
    .X(_01513_));
 sky130_fd_sc_hd__a22o_2 _15014_ (.A1(\core.instr_or ),
    .A2(_05932_),
    .B1(_05933_),
    .B2(_05945_),
    .X(_01941_));
 sky130_fd_sc_hd__and2_2 _15015_ (.A(_03546_),
    .B(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__buf_1 _15016_ (.A(_01942_),
    .X(_01514_));
 sky130_fd_sc_hd__a22o_2 _15017_ (.A1(\core.instr_srl ),
    .A2(_05932_),
    .B1(_05945_),
    .B2(_05953_),
    .X(_01943_));
 sky130_fd_sc_hd__and2_2 _15018_ (.A(_03546_),
    .B(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__buf_1 _15019_ (.A(_01944_),
    .X(_01515_));
 sky130_fd_sc_hd__a22o_2 _15020_ (.A1(\core.instr_sltu ),
    .A2(_05830_),
    .B1(_05929_),
    .B2(_05945_),
    .X(_01945_));
 sky130_fd_sc_hd__and2_2 _15021_ (.A(_03546_),
    .B(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__buf_1 _15022_ (.A(_01946_),
    .X(_01516_));
 sky130_fd_sc_hd__o2bb2a_2 _15023_ (.A1_N(\core.instr_slt ),
    .A2_N(_07089_),
    .B1(_05922_),
    .B2(_05948_),
    .X(_01947_));
 sky130_fd_sc_hd__nor2_2 _15024_ (.A(_02055_),
    .B(_01947_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_2 _15025_ (.A(_02912_),
    .B(_05877_),
    .Y(_01948_));
 sky130_fd_sc_hd__a41o_2 _15026_ (.A1(\core.mem_rdata_q[30] ),
    .A2(_05880_),
    .A3(_05940_),
    .A4(_05952_),
    .B1(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__and2_2 _15027_ (.A(_03546_),
    .B(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__buf_1 _15028_ (.A(_01950_),
    .X(_01518_));
 sky130_fd_sc_hd__a32o_2 _15029_ (.A1(_05878_),
    .A2(_05925_),
    .A3(_05942_),
    .B1(_05943_),
    .B2(\core.instr_slli ),
    .X(_01519_));
 sky130_fd_sc_hd__a22o_2 _15030_ (.A1(\core.instr_sw ),
    .A2(_05943_),
    .B1(_01931_),
    .B2(_02090_),
    .X(_01520_));
 sky130_fd_sc_hd__a22o_2 _15031_ (.A1(\core.instr_andi ),
    .A2(_05830_),
    .B1(_05925_),
    .B2(_01932_),
    .X(_01951_));
 sky130_fd_sc_hd__and2_2 _15032_ (.A(_03546_),
    .B(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__buf_1 _15033_ (.A(_01952_),
    .X(_01521_));
 sky130_fd_sc_hd__a32o_2 _15034_ (.A1(\core.mem_rdata_q[14] ),
    .A2(_05879_),
    .A3(_05925_),
    .B1(_05829_),
    .B2(\core.instr_xori ),
    .X(_01953_));
 sky130_fd_sc_hd__and2_2 _15035_ (.A(_03546_),
    .B(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__buf_1 _15036_ (.A(_01954_),
    .X(_01522_));
 sky130_fd_sc_hd__a22o_2 _15037_ (.A1(\core.instr_addi ),
    .A2(_05830_),
    .B1(_05880_),
    .B2(_05925_),
    .X(_01955_));
 sky130_fd_sc_hd__and2_2 _15038_ (.A(_03546_),
    .B(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__buf_1 _15039_ (.A(_01956_),
    .X(_01523_));
 sky130_fd_sc_hd__a22o_2 _15040_ (.A1(\core.instr_sb ),
    .A2(_05943_),
    .B1(_05881_),
    .B2(_02090_),
    .X(_01524_));
 sky130_fd_sc_hd__a22o_2 _15041_ (.A1(_02083_),
    .A2(_02051_),
    .B1(_05984_),
    .B2(\core.mem_do_rdata ),
    .X(_01525_));
 sky130_fd_sc_hd__and2_2 _15042_ (.A(_02236_),
    .B(_02445_),
    .X(_01957_));
 sky130_fd_sc_hd__inv_2 _15043_ (.A(_02091_),
    .Y(_01958_));
 sky130_fd_sc_hd__a31o_2 _15044_ (.A1(_01958_),
    .A2(\core.is_sll_srl_sra ),
    .A3(_02095_),
    .B1(_02092_),
    .X(_01959_));
 sky130_fd_sc_hd__a221oi_2 _15045_ (.A1(_02110_),
    .A2(_03471_),
    .B1(_01959_),
    .B2(\core.cpu_state[2] ),
    .C1(_02102_),
    .Y(_01960_));
 sky130_fd_sc_hd__nand2_2 _15046_ (.A(_02109_),
    .B(_03471_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21o_2 _15047_ (.A1(\core.is_sb_sh_sw ),
    .A2(_02094_),
    .B1(_02085_),
    .X(_01962_));
 sky130_fd_sc_hd__a211o_2 _15048_ (.A1(\core.cpu_state[2] ),
    .A2(_01962_),
    .B1(_03471_),
    .C1(\core.mem_do_prefetch ),
    .X(_01963_));
 sky130_fd_sc_hd__a21bo_2 _15049_ (.A1(_01961_),
    .A2(_01963_),
    .B1_N(_01960_),
    .X(_01964_));
 sky130_fd_sc_hd__o211a_2 _15050_ (.A1(\core.mem_do_rinst ),
    .A2(_01960_),
    .B1(_01964_),
    .C1(_05984_),
    .X(_01965_));
 sky130_fd_sc_hd__a31o_2 _15051_ (.A1(_01957_),
    .A2(_04424_),
    .A3(_05983_),
    .B1(_01965_),
    .X(_01526_));
 sky130_fd_sc_hd__inv_2 _15052_ (.A(\core.instr_jalr ),
    .Y(_01966_));
 sky130_fd_sc_hd__a21o_2 _15053_ (.A1(_02109_),
    .A2(_02111_),
    .B1(\core.mem_do_prefetch ),
    .X(_01967_));
 sky130_fd_sc_hd__o311a_2 _15054_ (.A1(_01966_),
    .A2(_03667_),
    .A3(_03791_),
    .B1(_05984_),
    .C1(_01967_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_2 _15055_ (.A0(\core.reg_out[2] ),
    .A1(\core.reg_next_pc[2] ),
    .S(_03245_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_2 _15056_ (.A0(_02372_),
    .A1(_01968_),
    .S(_03242_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_2 _15057_ (.A0(mem_addr[2]),
    .A1(_01969_),
    .S(_03236_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_1 _15058_ (.A(_01970_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_2 _15059_ (.A0(\core.reg_out[3] ),
    .A1(\core.reg_next_pc[3] ),
    .S(_03245_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_2 _15060_ (.A0(_02375_),
    .A1(_01971_),
    .S(_03242_),
    .X(_01972_));
 sky130_fd_sc_hd__buf_1 _15061_ (.A(_03213_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_2 _15062_ (.A0(mem_addr[3]),
    .A1(_01972_),
    .S(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__buf_1 _15063_ (.A(_01974_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_2 _15064_ (.A0(\core.reg_out[4] ),
    .A1(\core.reg_next_pc[4] ),
    .S(_03245_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_2 _15065_ (.A0(_02355_),
    .A1(_01975_),
    .S(_03242_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _15066_ (.A0(mem_addr[4]),
    .A1(_01976_),
    .S(_01973_),
    .X(_01977_));
 sky130_fd_sc_hd__buf_1 _15067_ (.A(_01977_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_2 _15068_ (.A0(\core.reg_out[5] ),
    .A1(\core.reg_next_pc[5] ),
    .S(_03245_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_2 _15069_ (.A0(_02388_),
    .A1(_01978_),
    .S(_03242_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_2 _15070_ (.A0(mem_addr[5]),
    .A1(_01979_),
    .S(_01973_),
    .X(_01980_));
 sky130_fd_sc_hd__buf_1 _15071_ (.A(_01980_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_2 _15072_ (.A0(\core.reg_out[6] ),
    .A1(\core.reg_next_pc[6] ),
    .S(_03245_),
    .X(_01981_));
 sky130_fd_sc_hd__buf_1 _15073_ (.A(_03206_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_2 _15074_ (.A0(_02383_),
    .A1(_01981_),
    .S(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_2 _15075_ (.A0(mem_addr[6]),
    .A1(_01983_),
    .S(_01973_),
    .X(_01984_));
 sky130_fd_sc_hd__buf_1 _15076_ (.A(_01984_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _15077_ (.A(_03202_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _15078_ (.A0(\core.reg_out[7] ),
    .A1(\core.reg_next_pc[7] ),
    .S(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_2 _15079_ (.A0(_02380_),
    .A1(_01986_),
    .S(_01982_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_2 _15080_ (.A0(mem_addr[7]),
    .A1(_01987_),
    .S(_01973_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_1 _15081_ (.A(_01988_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_2 _15082_ (.A0(\core.reg_out[8] ),
    .A1(\core.reg_next_pc[8] ),
    .S(_01985_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_2 _15083_ (.A0(_02327_),
    .A1(_01989_),
    .S(_01982_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_2 _15084_ (.A0(mem_addr[8]),
    .A1(_01990_),
    .S(_01973_),
    .X(_01991_));
 sky130_fd_sc_hd__buf_1 _15085_ (.A(_01991_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_2 _15086_ (.A0(\core.reg_out[9] ),
    .A1(\core.reg_next_pc[9] ),
    .S(_01985_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_2 _15087_ (.A0(_02331_),
    .A1(_01992_),
    .S(_01982_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_2 _15088_ (.A0(mem_addr[9]),
    .A1(_01993_),
    .S(_01973_),
    .X(_01994_));
 sky130_fd_sc_hd__buf_1 _15089_ (.A(_01994_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_2 _15090_ (.A0(\core.reg_out[10] ),
    .A1(\core.reg_next_pc[10] ),
    .S(_01985_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_2 _15091_ (.A0(_02323_),
    .A1(_01995_),
    .S(_01982_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_2 _15092_ (.A0(mem_addr[10]),
    .A1(_01996_),
    .S(_01973_),
    .X(_01997_));
 sky130_fd_sc_hd__buf_1 _15093_ (.A(_01997_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_2 _15094_ (.A0(\core.reg_out[11] ),
    .A1(\core.reg_next_pc[11] ),
    .S(_01985_),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_2 _15095_ (.A0(_02336_),
    .A1(_01998_),
    .S(_01982_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_2 _15096_ (.A0(mem_addr[11]),
    .A1(_01999_),
    .S(_01973_),
    .X(_02000_));
 sky130_fd_sc_hd__buf_1 _15097_ (.A(_02000_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_2 _15098_ (.A0(\core.reg_out[12] ),
    .A1(\core.reg_next_pc[12] ),
    .S(_01985_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_2 _15099_ (.A0(_02315_),
    .A1(_02001_),
    .S(_01982_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_2 _15100_ (.A0(mem_addr[12]),
    .A1(_02002_),
    .S(_01973_),
    .X(_02003_));
 sky130_fd_sc_hd__buf_1 _15101_ (.A(_02003_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_2 _15102_ (.A0(\core.reg_out[13] ),
    .A1(\core.reg_next_pc[13] ),
    .S(_01985_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_2 _15103_ (.A0(_02312_),
    .A1(_02004_),
    .S(_01982_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_2 _15104_ (.A0(mem_addr[13]),
    .A1(_02005_),
    .S(_03213_),
    .X(_02006_));
 sky130_fd_sc_hd__buf_1 _15105_ (.A(_02006_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_2 _15106_ (.A0(\core.reg_out[14] ),
    .A1(\core.reg_next_pc[14] ),
    .S(_01985_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_2 _15107_ (.A0(_02306_),
    .A1(_02007_),
    .S(_01982_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_2 _15108_ (.A0(mem_addr[14]),
    .A1(_02008_),
    .S(_03213_),
    .X(_02009_));
 sky130_fd_sc_hd__buf_1 _15109_ (.A(_02009_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_2 _15110_ (.A0(\core.reg_out[15] ),
    .A1(\core.reg_next_pc[15] ),
    .S(_01985_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_2 _15111_ (.A0(_02345_),
    .A1(_02010_),
    .S(_01982_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_2 _15112_ (.A0(mem_addr[15]),
    .A1(_02011_),
    .S(_03213_),
    .X(_02012_));
 sky130_fd_sc_hd__buf_1 _15113_ (.A(_02012_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_2 _15114_ (.A0(\core.reg_out[16] ),
    .A1(\core.reg_next_pc[16] ),
    .S(_01985_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_2 _15115_ (.A0(_02291_),
    .A1(_02013_),
    .S(_03206_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_2 _15116_ (.A0(mem_addr[16]),
    .A1(_02014_),
    .S(_03213_),
    .X(_02015_));
 sky130_fd_sc_hd__buf_1 _15117_ (.A(_02015_),
    .X(_01542_));
 sky130_fd_sc_hd__dfxtp_2 _15118_ (.CLK(clk),
    .D(_00037_),
    .Q(mem_addr[17]));
 sky130_fd_sc_hd__dfxtp_2 _15119_ (.CLK(clk),
    .D(_00038_),
    .Q(mem_addr[18]));
 sky130_fd_sc_hd__dfxtp_2 _15120_ (.CLK(clk),
    .D(_00039_),
    .Q(mem_addr[19]));
 sky130_fd_sc_hd__dfxtp_2 _15121_ (.CLK(clk),
    .D(_00040_),
    .Q(mem_addr[20]));
 sky130_fd_sc_hd__dfxtp_2 _15122_ (.CLK(clk),
    .D(_00041_),
    .Q(mem_addr[21]));
 sky130_fd_sc_hd__dfxtp_2 _15123_ (.CLK(clk),
    .D(_00042_),
    .Q(mem_addr[22]));
 sky130_fd_sc_hd__dfxtp_2 _15124_ (.CLK(clk),
    .D(_00043_),
    .Q(mem_addr[23]));
 sky130_fd_sc_hd__dfxtp_2 _15125_ (.CLK(clk),
    .D(_00044_),
    .Q(mem_addr[24]));
 sky130_fd_sc_hd__dfxtp_2 _15126_ (.CLK(clk),
    .D(_00045_),
    .Q(mem_addr[25]));
 sky130_fd_sc_hd__dfxtp_2 _15127_ (.CLK(clk),
    .D(_00046_),
    .Q(mem_addr[26]));
 sky130_fd_sc_hd__dfxtp_2 _15128_ (.CLK(clk),
    .D(_00047_),
    .Q(mem_addr[27]));
 sky130_fd_sc_hd__dfxtp_2 _15129_ (.CLK(clk),
    .D(_00048_),
    .Q(mem_addr[28]));
 sky130_fd_sc_hd__dfxtp_2 _15130_ (.CLK(clk),
    .D(_00049_),
    .Q(mem_addr[29]));
 sky130_fd_sc_hd__dfxtp_2 _15131_ (.CLK(clk),
    .D(_00050_),
    .Q(mem_addr[30]));
 sky130_fd_sc_hd__dfxtp_2 _15132_ (.CLK(clk),
    .D(_00051_),
    .Q(mem_addr[31]));
 sky130_fd_sc_hd__dfxtp_2 _15133_ (.CLK(clk),
    .D(_01543_),
    .Q(\core.reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15134_ (.CLK(clk),
    .D(_01554_),
    .Q(\core.reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15135_ (.CLK(clk),
    .D(_01565_),
    .Q(\core.reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15136_ (.CLK(clk),
    .D(_01568_),
    .Q(\core.reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15137_ (.CLK(clk),
    .D(_01569_),
    .Q(\core.reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15138_ (.CLK(clk),
    .D(_01570_),
    .Q(\core.reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15139_ (.CLK(clk),
    .D(_01571_),
    .Q(\core.reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15140_ (.CLK(clk),
    .D(_01572_),
    .Q(\core.reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15141_ (.CLK(clk),
    .D(_01573_),
    .Q(\core.reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15142_ (.CLK(clk),
    .D(_01574_),
    .Q(\core.reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15143_ (.CLK(clk),
    .D(_01544_),
    .Q(\core.reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15144_ (.CLK(clk),
    .D(_01545_),
    .Q(\core.reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15145_ (.CLK(clk),
    .D(_01546_),
    .Q(\core.reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15146_ (.CLK(clk),
    .D(_01547_),
    .Q(\core.reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15147_ (.CLK(clk),
    .D(_01548_),
    .Q(\core.reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15148_ (.CLK(clk),
    .D(_01549_),
    .Q(\core.reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15149_ (.CLK(clk),
    .D(_01550_),
    .Q(\core.reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15150_ (.CLK(clk),
    .D(_01551_),
    .Q(\core.reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15151_ (.CLK(clk),
    .D(_01552_),
    .Q(\core.reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15152_ (.CLK(clk),
    .D(_01553_),
    .Q(\core.reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15153_ (.CLK(clk),
    .D(_01555_),
    .Q(\core.reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15154_ (.CLK(clk),
    .D(_01556_),
    .Q(\core.reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15155_ (.CLK(clk),
    .D(_01557_),
    .Q(\core.reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15156_ (.CLK(clk),
    .D(_01558_),
    .Q(\core.reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15157_ (.CLK(clk),
    .D(_01559_),
    .Q(\core.reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15158_ (.CLK(clk),
    .D(_01560_),
    .Q(\core.reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15159_ (.CLK(clk),
    .D(_01561_),
    .Q(\core.reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15160_ (.CLK(clk),
    .D(_01562_),
    .Q(\core.reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15161_ (.CLK(clk),
    .D(_01563_),
    .Q(\core.reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15162_ (.CLK(clk),
    .D(_01564_),
    .Q(\core.reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15163_ (.CLK(clk),
    .D(_01566_),
    .Q(\core.reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15164_ (.CLK(clk),
    .D(_01567_),
    .Q(\core.reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15165_ (.CLK(clk),
    .D(_00052_),
    .Q(\core.pcpi_rs1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15166_ (.CLK(clk),
    .D(_00053_),
    .Q(\core.count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15167_ (.CLK(clk),
    .D(_00054_),
    .Q(\core.count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15168_ (.CLK(clk),
    .D(_00055_),
    .Q(\core.count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15169_ (.CLK(clk),
    .D(_00056_),
    .Q(\core.count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15170_ (.CLK(clk),
    .D(_00057_),
    .Q(\core.count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15171_ (.CLK(clk),
    .D(_00058_),
    .Q(\core.count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15172_ (.CLK(clk),
    .D(_00059_),
    .Q(\core.count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15173_ (.CLK(clk),
    .D(_00060_),
    .Q(\core.count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15174_ (.CLK(clk),
    .D(_00061_),
    .Q(\core.count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15175_ (.CLK(clk),
    .D(_00062_),
    .Q(\core.count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15176_ (.CLK(clk),
    .D(_00063_),
    .Q(\core.count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15177_ (.CLK(clk),
    .D(_00064_),
    .Q(\core.count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15178_ (.CLK(clk),
    .D(_00065_),
    .Q(\core.count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15179_ (.CLK(clk),
    .D(_00066_),
    .Q(\core.count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15180_ (.CLK(clk),
    .D(_00067_),
    .Q(\core.count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15181_ (.CLK(clk),
    .D(_00068_),
    .Q(\core.count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15182_ (.CLK(clk),
    .D(_00069_),
    .Q(\core.count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15183_ (.CLK(clk),
    .D(_00070_),
    .Q(\core.count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15184_ (.CLK(clk),
    .D(_00071_),
    .Q(\core.count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15185_ (.CLK(clk),
    .D(_00072_),
    .Q(\core.count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15186_ (.CLK(clk),
    .D(_00073_),
    .Q(\core.count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15187_ (.CLK(clk),
    .D(_00074_),
    .Q(\core.count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15188_ (.CLK(clk),
    .D(_00075_),
    .Q(\core.count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15189_ (.CLK(clk),
    .D(_00076_),
    .Q(\core.count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15190_ (.CLK(clk),
    .D(_00077_),
    .Q(\core.count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15191_ (.CLK(clk),
    .D(_00078_),
    .Q(\core.count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15192_ (.CLK(clk),
    .D(_00079_),
    .Q(\core.count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15193_ (.CLK(clk),
    .D(_00080_),
    .Q(\core.count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15194_ (.CLK(clk),
    .D(_00081_),
    .Q(\core.count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15195_ (.CLK(clk),
    .D(_00082_),
    .Q(\core.count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15196_ (.CLK(clk),
    .D(_00083_),
    .Q(\core.count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15197_ (.CLK(clk),
    .D(_00084_),
    .Q(\core.count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15198_ (.CLK(clk),
    .D(_00085_),
    .Q(\core.count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_2 _15199_ (.CLK(clk),
    .D(_00086_),
    .Q(\core.count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_2 _15200_ (.CLK(clk),
    .D(_00087_),
    .Q(\core.count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_2 _15201_ (.CLK(clk),
    .D(_00088_),
    .Q(\core.count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_2 _15202_ (.CLK(clk),
    .D(_00089_),
    .Q(\core.count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_2 _15203_ (.CLK(clk),
    .D(_00090_),
    .Q(\core.count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_2 _15204_ (.CLK(clk),
    .D(_00091_),
    .Q(\core.count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_2 _15205_ (.CLK(clk),
    .D(_00092_),
    .Q(\core.count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_2 _15206_ (.CLK(clk),
    .D(_00093_),
    .Q(\core.count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_2 _15207_ (.CLK(clk),
    .D(_00094_),
    .Q(\core.count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_2 _15208_ (.CLK(clk),
    .D(_00095_),
    .Q(\core.count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_2 _15209_ (.CLK(clk),
    .D(_00096_),
    .Q(\core.count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_2 _15210_ (.CLK(clk),
    .D(_00097_),
    .Q(\core.count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_2 _15211_ (.CLK(clk),
    .D(_00098_),
    .Q(\core.count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_2 _15212_ (.CLK(clk),
    .D(_00099_),
    .Q(\core.count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_2 _15213_ (.CLK(clk),
    .D(_00100_),
    .Q(\core.count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_2 _15214_ (.CLK(clk),
    .D(_00101_),
    .Q(\core.count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_2 _15215_ (.CLK(clk),
    .D(_00102_),
    .Q(\core.count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_2 _15216_ (.CLK(clk),
    .D(_00103_),
    .Q(\core.count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_2 _15217_ (.CLK(clk),
    .D(_00104_),
    .Q(\core.count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_2 _15218_ (.CLK(clk),
    .D(_00105_),
    .Q(\core.count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 _15219_ (.CLK(clk),
    .D(_00106_),
    .Q(\core.count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_2 _15220_ (.CLK(clk),
    .D(_00107_),
    .Q(\core.count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_2 _15221_ (.CLK(clk),
    .D(_00108_),
    .Q(\core.count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_2 _15222_ (.CLK(clk),
    .D(_00109_),
    .Q(\core.count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_2 _15223_ (.CLK(clk),
    .D(_00110_),
    .Q(\core.count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_2 _15224_ (.CLK(clk),
    .D(_00111_),
    .Q(\core.count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_2 _15225_ (.CLK(clk),
    .D(_00112_),
    .Q(\core.count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_2 _15226_ (.CLK(clk),
    .D(_00113_),
    .Q(\core.count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_2 _15227_ (.CLK(clk),
    .D(_00114_),
    .Q(\core.count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_2 _15228_ (.CLK(clk),
    .D(_00115_),
    .Q(\core.count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_2 _15229_ (.CLK(clk),
    .D(_00116_),
    .Q(\core.count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_2 _15230_ (.CLK(clk),
    .D(_00117_),
    .Q(\core.reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15231_ (.CLK(clk),
    .D(_00118_),
    .Q(\core.reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15232_ (.CLK(clk),
    .D(_00119_),
    .Q(\core.reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15233_ (.CLK(clk),
    .D(_00120_),
    .Q(\core.reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15234_ (.CLK(clk),
    .D(_00121_),
    .Q(\core.reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15235_ (.CLK(clk),
    .D(_00122_),
    .Q(\core.reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15236_ (.CLK(clk),
    .D(_00123_),
    .Q(\core.reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15237_ (.CLK(clk),
    .D(_00124_),
    .Q(\core.reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15238_ (.CLK(clk),
    .D(_00125_),
    .Q(\core.reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15239_ (.CLK(clk),
    .D(_00126_),
    .Q(\core.reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15240_ (.CLK(clk),
    .D(_00127_),
    .Q(\core.reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15241_ (.CLK(clk),
    .D(_00128_),
    .Q(\core.reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15242_ (.CLK(clk),
    .D(_00129_),
    .Q(\core.reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15243_ (.CLK(clk),
    .D(_00130_),
    .Q(\core.reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15244_ (.CLK(clk),
    .D(_00131_),
    .Q(\core.reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15245_ (.CLK(clk),
    .D(_00132_),
    .Q(\core.reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15246_ (.CLK(clk),
    .D(_00133_),
    .Q(\core.reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15247_ (.CLK(clk),
    .D(_00134_),
    .Q(\core.reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15248_ (.CLK(clk),
    .D(_00135_),
    .Q(\core.reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15249_ (.CLK(clk),
    .D(_00136_),
    .Q(\core.reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15250_ (.CLK(clk),
    .D(_00137_),
    .Q(\core.reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15251_ (.CLK(clk),
    .D(_00138_),
    .Q(\core.reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15252_ (.CLK(clk),
    .D(_00139_),
    .Q(\core.reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15253_ (.CLK(clk),
    .D(_00140_),
    .Q(\core.reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15254_ (.CLK(clk),
    .D(_00141_),
    .Q(\core.reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15255_ (.CLK(clk),
    .D(_00142_),
    .Q(\core.reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15256_ (.CLK(clk),
    .D(_00143_),
    .Q(\core.reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15257_ (.CLK(clk),
    .D(_00144_),
    .Q(\core.reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15258_ (.CLK(clk),
    .D(_00145_),
    .Q(\core.reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15259_ (.CLK(clk),
    .D(_00146_),
    .Q(\core.reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15260_ (.CLK(clk),
    .D(_00147_),
    .Q(\core.reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15261_ (.CLK(clk),
    .D(_00148_),
    .Q(\core.reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15262_ (.CLK(clk),
    .D(_00149_),
    .Q(\core.reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15263_ (.CLK(clk),
    .D(_00150_),
    .Q(\core.reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15264_ (.CLK(clk),
    .D(_00151_),
    .Q(\core.reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15265_ (.CLK(clk),
    .D(_00152_),
    .Q(\core.reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15266_ (.CLK(clk),
    .D(_00153_),
    .Q(\core.reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15267_ (.CLK(clk),
    .D(_00154_),
    .Q(\core.reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15268_ (.CLK(clk),
    .D(_00155_),
    .Q(\core.reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15269_ (.CLK(clk),
    .D(_00156_),
    .Q(\core.reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15270_ (.CLK(clk),
    .D(_00157_),
    .Q(\core.reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15271_ (.CLK(clk),
    .D(_00158_),
    .Q(\core.reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15272_ (.CLK(clk),
    .D(_00159_),
    .Q(\core.reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15273_ (.CLK(clk),
    .D(_00160_),
    .Q(\core.reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15274_ (.CLK(clk),
    .D(_00161_),
    .Q(\core.reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15275_ (.CLK(clk),
    .D(_00162_),
    .Q(\core.reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15276_ (.CLK(clk),
    .D(_00163_),
    .Q(\core.reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15277_ (.CLK(clk),
    .D(_00164_),
    .Q(\core.reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15278_ (.CLK(clk),
    .D(_00165_),
    .Q(\core.reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15279_ (.CLK(clk),
    .D(_00166_),
    .Q(\core.reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15280_ (.CLK(clk),
    .D(_00167_),
    .Q(\core.reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15281_ (.CLK(clk),
    .D(_00168_),
    .Q(\core.reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15282_ (.CLK(clk),
    .D(_00169_),
    .Q(\core.reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15283_ (.CLK(clk),
    .D(_00170_),
    .Q(\core.reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15284_ (.CLK(clk),
    .D(_00171_),
    .Q(\core.reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15285_ (.CLK(clk),
    .D(_00172_),
    .Q(\core.reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15286_ (.CLK(clk),
    .D(_00173_),
    .Q(\core.reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15287_ (.CLK(clk),
    .D(_00174_),
    .Q(\core.reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15288_ (.CLK(clk),
    .D(_00175_),
    .Q(\core.reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15289_ (.CLK(clk),
    .D(_00176_),
    .Q(\core.reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15290_ (.CLK(clk),
    .D(_00177_),
    .Q(\core.reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15291_ (.CLK(clk),
    .D(_00178_),
    .Q(\core.reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15292_ (.CLK(clk),
    .D(_00179_),
    .Q(\core.count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15293_ (.CLK(clk),
    .D(_00180_),
    .Q(\core.count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15294_ (.CLK(clk),
    .D(_00181_),
    .Q(\core.count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15295_ (.CLK(clk),
    .D(_00182_),
    .Q(\core.count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15296_ (.CLK(clk),
    .D(_00183_),
    .Q(\core.count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15297_ (.CLK(clk),
    .D(_00184_),
    .Q(\core.count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15298_ (.CLK(clk),
    .D(_00185_),
    .Q(\core.count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15299_ (.CLK(clk),
    .D(_00186_),
    .Q(\core.count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15300_ (.CLK(clk),
    .D(_00187_),
    .Q(\core.count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15301_ (.CLK(clk),
    .D(_00188_),
    .Q(\core.count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15302_ (.CLK(clk),
    .D(_00189_),
    .Q(\core.count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15303_ (.CLK(clk),
    .D(_00190_),
    .Q(\core.count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15304_ (.CLK(clk),
    .D(_00191_),
    .Q(\core.count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15305_ (.CLK(clk),
    .D(_00192_),
    .Q(\core.count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15306_ (.CLK(clk),
    .D(_00193_),
    .Q(\core.count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15307_ (.CLK(clk),
    .D(_00194_),
    .Q(\core.count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15308_ (.CLK(clk),
    .D(_00195_),
    .Q(\core.count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15309_ (.CLK(clk),
    .D(_00196_),
    .Q(\core.count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15310_ (.CLK(clk),
    .D(_00197_),
    .Q(\core.count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15311_ (.CLK(clk),
    .D(_00198_),
    .Q(\core.count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15312_ (.CLK(clk),
    .D(_00199_),
    .Q(\core.count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15313_ (.CLK(clk),
    .D(_00200_),
    .Q(\core.count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15314_ (.CLK(clk),
    .D(_00201_),
    .Q(\core.count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15315_ (.CLK(clk),
    .D(_00202_),
    .Q(\core.count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15316_ (.CLK(clk),
    .D(_00203_),
    .Q(\core.count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15317_ (.CLK(clk),
    .D(_00204_),
    .Q(\core.count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15318_ (.CLK(clk),
    .D(_00205_),
    .Q(\core.count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15319_ (.CLK(clk),
    .D(_00206_),
    .Q(\core.count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15320_ (.CLK(clk),
    .D(_00207_),
    .Q(\core.count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15321_ (.CLK(clk),
    .D(_00208_),
    .Q(\core.count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15322_ (.CLK(clk),
    .D(_00209_),
    .Q(\core.count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15323_ (.CLK(clk),
    .D(_00210_),
    .Q(\core.count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15324_ (.CLK(clk),
    .D(_00211_),
    .Q(\core.count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_2 _15325_ (.CLK(clk),
    .D(_00212_),
    .Q(\core.count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_2 _15326_ (.CLK(clk),
    .D(_00213_),
    .Q(\core.count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_2 _15327_ (.CLK(clk),
    .D(_00214_),
    .Q(\core.count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_2 _15328_ (.CLK(clk),
    .D(_00215_),
    .Q(\core.count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_2 _15329_ (.CLK(clk),
    .D(_00216_),
    .Q(\core.count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_2 _15330_ (.CLK(clk),
    .D(_00217_),
    .Q(\core.count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_2 _15331_ (.CLK(clk),
    .D(_00218_),
    .Q(\core.count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_2 _15332_ (.CLK(clk),
    .D(_00219_),
    .Q(\core.count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_2 _15333_ (.CLK(clk),
    .D(_00220_),
    .Q(\core.count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_2 _15334_ (.CLK(clk),
    .D(_00221_),
    .Q(\core.count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_2 _15335_ (.CLK(clk),
    .D(_00222_),
    .Q(\core.count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_2 _15336_ (.CLK(clk),
    .D(_00223_),
    .Q(\core.count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_2 _15337_ (.CLK(clk),
    .D(_00224_),
    .Q(\core.count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_2 _15338_ (.CLK(clk),
    .D(_00225_),
    .Q(\core.count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_2 _15339_ (.CLK(clk),
    .D(_00226_),
    .Q(\core.count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_2 _15340_ (.CLK(clk),
    .D(_00227_),
    .Q(\core.count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_2 _15341_ (.CLK(clk),
    .D(_00228_),
    .Q(\core.count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_2 _15342_ (.CLK(clk),
    .D(_00229_),
    .Q(\core.count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_2 _15343_ (.CLK(clk),
    .D(_00230_),
    .Q(\core.count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_2 _15344_ (.CLK(clk),
    .D(_00231_),
    .Q(\core.count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_2 _15345_ (.CLK(clk),
    .D(_00232_),
    .Q(\core.count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_2 _15346_ (.CLK(clk),
    .D(_00233_),
    .Q(\core.count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_2 _15347_ (.CLK(clk),
    .D(_00234_),
    .Q(\core.count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_2 _15348_ (.CLK(clk),
    .D(_00235_),
    .Q(\core.count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_2 _15349_ (.CLK(clk),
    .D(_00236_),
    .Q(\core.count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_2 _15350_ (.CLK(clk),
    .D(_00237_),
    .Q(\core.count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_2 _15351_ (.CLK(clk),
    .D(_00238_),
    .Q(\core.count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_2 _15352_ (.CLK(clk),
    .D(_00239_),
    .Q(\core.count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_2 _15353_ (.CLK(clk),
    .D(_00240_),
    .Q(\core.count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_2 _15354_ (.CLK(clk),
    .D(_00241_),
    .Q(\core.count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_2 _15355_ (.CLK(clk),
    .D(_00242_),
    .Q(\core.count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_2 _15356_ (.CLK(clk),
    .D(_00243_),
    .Q(\core.pcpi_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15357_ (.CLK(clk),
    .D(_00244_),
    .Q(\core.pcpi_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15358_ (.CLK(clk),
    .D(_00245_),
    .Q(\core.pcpi_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15359_ (.CLK(clk),
    .D(_00246_),
    .Q(\core.pcpi_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15360_ (.CLK(clk),
    .D(_00247_),
    .Q(\core.pcpi_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15361_ (.CLK(clk),
    .D(_00248_),
    .Q(\core.pcpi_rs1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15362_ (.CLK(clk),
    .D(_00249_),
    .Q(\core.pcpi_rs1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15363_ (.CLK(clk),
    .D(_00250_),
    .Q(\core.pcpi_rs1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15364_ (.CLK(clk),
    .D(_00251_),
    .Q(\core.pcpi_rs1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15365_ (.CLK(clk),
    .D(_00252_),
    .Q(\core.pcpi_rs1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15366_ (.CLK(clk),
    .D(_00253_),
    .Q(\core.pcpi_rs1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15367_ (.CLK(clk),
    .D(_00254_),
    .Q(\core.pcpi_rs1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15368_ (.CLK(clk),
    .D(_00255_),
    .Q(\core.pcpi_rs1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15369_ (.CLK(clk),
    .D(_00256_),
    .Q(\core.pcpi_rs1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15370_ (.CLK(clk),
    .D(_00257_),
    .Q(\core.pcpi_rs1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15371_ (.CLK(clk),
    .D(_00258_),
    .Q(\core.pcpi_rs1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15372_ (.CLK(clk),
    .D(_00259_),
    .Q(\core.pcpi_rs1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15373_ (.CLK(clk),
    .D(_00260_),
    .Q(\core.pcpi_rs1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15374_ (.CLK(clk),
    .D(_00261_),
    .Q(\core.pcpi_rs1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15375_ (.CLK(clk),
    .D(_00262_),
    .Q(\core.pcpi_rs1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15376_ (.CLK(clk),
    .D(_00263_),
    .Q(\core.pcpi_rs1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15377_ (.CLK(clk),
    .D(_00264_),
    .Q(\core.pcpi_rs1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15378_ (.CLK(clk),
    .D(_00265_),
    .Q(\core.pcpi_rs1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15379_ (.CLK(clk),
    .D(_00266_),
    .Q(\core.pcpi_rs1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15380_ (.CLK(clk),
    .D(_00267_),
    .Q(\core.pcpi_rs1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15381_ (.CLK(clk),
    .D(_00268_),
    .Q(\core.pcpi_rs1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15382_ (.CLK(clk),
    .D(_00269_),
    .Q(\core.pcpi_rs1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15383_ (.CLK(clk),
    .D(_00270_),
    .Q(\core.pcpi_rs1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15384_ (.CLK(clk),
    .D(_00271_),
    .Q(\core.pcpi_rs1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15385_ (.CLK(clk),
    .D(_00272_),
    .Q(\core.pcpi_rs1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15386_ (.CLK(clk),
    .D(_00273_),
    .Q(\core.pcpi_rs1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15387_ (.CLK(clk),
    .D(_00274_),
    .Q(\core.mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15388_ (.CLK(clk),
    .D(_00275_),
    .Q(\core.mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15389_ (.CLK(clk),
    .D(_00276_),
    .Q(\core.cpuregs[23][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15390_ (.CLK(clk),
    .D(_00277_),
    .Q(\core.cpuregs[23][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15391_ (.CLK(clk),
    .D(_00278_),
    .Q(\core.cpuregs[23][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15392_ (.CLK(clk),
    .D(_00279_),
    .Q(\core.cpuregs[23][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15393_ (.CLK(clk),
    .D(_00280_),
    .Q(\core.cpuregs[23][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15394_ (.CLK(clk),
    .D(_00281_),
    .Q(\core.cpuregs[23][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15395_ (.CLK(clk),
    .D(_00282_),
    .Q(\core.cpuregs[23][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15396_ (.CLK(clk),
    .D(_00283_),
    .Q(\core.cpuregs[23][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15397_ (.CLK(clk),
    .D(_00284_),
    .Q(\core.cpuregs[23][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15398_ (.CLK(clk),
    .D(_00285_),
    .Q(\core.cpuregs[23][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15399_ (.CLK(clk),
    .D(_00286_),
    .Q(\core.cpuregs[23][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15400_ (.CLK(clk),
    .D(_00287_),
    .Q(\core.cpuregs[23][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15401_ (.CLK(clk),
    .D(_00288_),
    .Q(\core.cpuregs[23][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15402_ (.CLK(clk),
    .D(_00289_),
    .Q(\core.cpuregs[23][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15403_ (.CLK(clk),
    .D(_00290_),
    .Q(\core.cpuregs[23][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15404_ (.CLK(clk),
    .D(_00291_),
    .Q(\core.cpuregs[23][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15405_ (.CLK(clk),
    .D(_00292_),
    .Q(\core.cpuregs[23][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15406_ (.CLK(clk),
    .D(_00293_),
    .Q(\core.cpuregs[23][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15407_ (.CLK(clk),
    .D(_00294_),
    .Q(\core.cpuregs[23][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15408_ (.CLK(clk),
    .D(_00295_),
    .Q(\core.cpuregs[23][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15409_ (.CLK(clk),
    .D(_00296_),
    .Q(\core.cpuregs[23][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15410_ (.CLK(clk),
    .D(_00297_),
    .Q(\core.cpuregs[23][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15411_ (.CLK(clk),
    .D(_00298_),
    .Q(\core.cpuregs[23][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15412_ (.CLK(clk),
    .D(_00299_),
    .Q(\core.cpuregs[23][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15413_ (.CLK(clk),
    .D(_00300_),
    .Q(\core.cpuregs[23][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15414_ (.CLK(clk),
    .D(_00301_),
    .Q(\core.cpuregs[23][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15415_ (.CLK(clk),
    .D(_00302_),
    .Q(\core.cpuregs[23][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15416_ (.CLK(clk),
    .D(_00303_),
    .Q(\core.cpuregs[23][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15417_ (.CLK(clk),
    .D(_00304_),
    .Q(\core.cpuregs[23][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15418_ (.CLK(clk),
    .D(_00305_),
    .Q(\core.cpuregs[23][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15419_ (.CLK(clk),
    .D(_00306_),
    .Q(\core.cpuregs[23][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15420_ (.CLK(clk),
    .D(_00307_),
    .Q(\core.cpuregs[23][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15421_ (.CLK(clk),
    .D(_00308_),
    .Q(\core.cpuregs[30][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15422_ (.CLK(clk),
    .D(_00309_),
    .Q(\core.cpuregs[30][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15423_ (.CLK(clk),
    .D(_00310_),
    .Q(\core.cpuregs[30][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15424_ (.CLK(clk),
    .D(_00311_),
    .Q(\core.cpuregs[30][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15425_ (.CLK(clk),
    .D(_00312_),
    .Q(\core.cpuregs[30][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15426_ (.CLK(clk),
    .D(_00313_),
    .Q(\core.cpuregs[30][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15427_ (.CLK(clk),
    .D(_00314_),
    .Q(\core.cpuregs[30][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15428_ (.CLK(clk),
    .D(_00315_),
    .Q(\core.cpuregs[30][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15429_ (.CLK(clk),
    .D(_00316_),
    .Q(\core.cpuregs[30][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15430_ (.CLK(clk),
    .D(_00317_),
    .Q(\core.cpuregs[30][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15431_ (.CLK(clk),
    .D(_00318_),
    .Q(\core.cpuregs[30][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15432_ (.CLK(clk),
    .D(_00319_),
    .Q(\core.cpuregs[30][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15433_ (.CLK(clk),
    .D(_00320_),
    .Q(\core.cpuregs[30][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15434_ (.CLK(clk),
    .D(_00321_),
    .Q(\core.cpuregs[30][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15435_ (.CLK(clk),
    .D(_00322_),
    .Q(\core.cpuregs[30][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15436_ (.CLK(clk),
    .D(_00323_),
    .Q(\core.cpuregs[30][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15437_ (.CLK(clk),
    .D(_00324_),
    .Q(\core.cpuregs[30][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15438_ (.CLK(clk),
    .D(_00325_),
    .Q(\core.cpuregs[30][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15439_ (.CLK(clk),
    .D(_00326_),
    .Q(\core.cpuregs[30][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15440_ (.CLK(clk),
    .D(_00327_),
    .Q(\core.cpuregs[30][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15441_ (.CLK(clk),
    .D(_00328_),
    .Q(\core.cpuregs[30][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15442_ (.CLK(clk),
    .D(_00329_),
    .Q(\core.cpuregs[30][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15443_ (.CLK(clk),
    .D(_00330_),
    .Q(\core.cpuregs[30][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15444_ (.CLK(clk),
    .D(_00331_),
    .Q(\core.cpuregs[30][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15445_ (.CLK(clk),
    .D(_00332_),
    .Q(\core.cpuregs[30][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15446_ (.CLK(clk),
    .D(_00333_),
    .Q(\core.cpuregs[30][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15447_ (.CLK(clk),
    .D(_00334_),
    .Q(\core.cpuregs[30][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15448_ (.CLK(clk),
    .D(_00335_),
    .Q(\core.cpuregs[30][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15449_ (.CLK(clk),
    .D(_00336_),
    .Q(\core.cpuregs[30][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15450_ (.CLK(clk),
    .D(_00337_),
    .Q(\core.cpuregs[30][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15451_ (.CLK(clk),
    .D(_00338_),
    .Q(\core.cpuregs[30][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15452_ (.CLK(clk),
    .D(_00339_),
    .Q(\core.cpuregs[30][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15453_ (.CLK(clk),
    .D(_00340_),
    .Q(\core.reg_sh[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15454_ (.CLK(clk),
    .D(_00341_),
    .Q(\core.reg_sh[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15455_ (.CLK(clk),
    .D(_00342_),
    .Q(\core.cpuregs[22][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15456_ (.CLK(clk),
    .D(_00343_),
    .Q(\core.cpuregs[22][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15457_ (.CLK(clk),
    .D(_00344_),
    .Q(\core.cpuregs[22][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15458_ (.CLK(clk),
    .D(_00345_),
    .Q(\core.cpuregs[22][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15459_ (.CLK(clk),
    .D(_00346_),
    .Q(\core.cpuregs[22][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15460_ (.CLK(clk),
    .D(_00347_),
    .Q(\core.cpuregs[22][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15461_ (.CLK(clk),
    .D(_00348_),
    .Q(\core.cpuregs[22][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15462_ (.CLK(clk),
    .D(_00349_),
    .Q(\core.cpuregs[22][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15463_ (.CLK(clk),
    .D(_00350_),
    .Q(\core.cpuregs[22][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15464_ (.CLK(clk),
    .D(_00351_),
    .Q(\core.cpuregs[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15465_ (.CLK(clk),
    .D(_00352_),
    .Q(\core.cpuregs[22][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15466_ (.CLK(clk),
    .D(_00353_),
    .Q(\core.cpuregs[22][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15467_ (.CLK(clk),
    .D(_00354_),
    .Q(\core.cpuregs[22][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15468_ (.CLK(clk),
    .D(_00355_),
    .Q(\core.cpuregs[22][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15469_ (.CLK(clk),
    .D(_00356_),
    .Q(\core.cpuregs[22][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15470_ (.CLK(clk),
    .D(_00357_),
    .Q(\core.cpuregs[22][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15471_ (.CLK(clk),
    .D(_00358_),
    .Q(\core.cpuregs[22][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15472_ (.CLK(clk),
    .D(_00359_),
    .Q(\core.cpuregs[22][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15473_ (.CLK(clk),
    .D(_00360_),
    .Q(\core.cpuregs[22][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15474_ (.CLK(clk),
    .D(_00361_),
    .Q(\core.cpuregs[22][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15475_ (.CLK(clk),
    .D(_00362_),
    .Q(\core.cpuregs[22][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15476_ (.CLK(clk),
    .D(_00363_),
    .Q(\core.cpuregs[22][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15477_ (.CLK(clk),
    .D(_00364_),
    .Q(\core.cpuregs[22][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15478_ (.CLK(clk),
    .D(_00365_),
    .Q(\core.cpuregs[22][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15479_ (.CLK(clk),
    .D(_00366_),
    .Q(\core.cpuregs[22][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15480_ (.CLK(clk),
    .D(_00367_),
    .Q(\core.cpuregs[22][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15481_ (.CLK(clk),
    .D(_00368_),
    .Q(\core.cpuregs[22][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15482_ (.CLK(clk),
    .D(_00369_),
    .Q(\core.cpuregs[22][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15483_ (.CLK(clk),
    .D(_00370_),
    .Q(\core.cpuregs[22][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15484_ (.CLK(clk),
    .D(_00371_),
    .Q(\core.cpuregs[22][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15485_ (.CLK(clk),
    .D(_00372_),
    .Q(\core.cpuregs[22][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15486_ (.CLK(clk),
    .D(_00373_),
    .Q(\core.cpuregs[22][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15487_ (.CLK(clk),
    .D(_00374_),
    .Q(\core.cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15488_ (.CLK(clk),
    .D(_00375_),
    .Q(\core.cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15489_ (.CLK(clk),
    .D(_00376_),
    .Q(\core.cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15490_ (.CLK(clk),
    .D(_00377_),
    .Q(\core.cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15491_ (.CLK(clk),
    .D(_00378_),
    .Q(\core.cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15492_ (.CLK(clk),
    .D(_00379_),
    .Q(\core.cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15493_ (.CLK(clk),
    .D(_00380_),
    .Q(\core.cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15494_ (.CLK(clk),
    .D(_00381_),
    .Q(\core.cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15495_ (.CLK(clk),
    .D(_00382_),
    .Q(\core.cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15496_ (.CLK(clk),
    .D(_00383_),
    .Q(\core.cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15497_ (.CLK(clk),
    .D(_00384_),
    .Q(\core.cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15498_ (.CLK(clk),
    .D(_00385_),
    .Q(\core.cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15499_ (.CLK(clk),
    .D(_00386_),
    .Q(\core.cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15500_ (.CLK(clk),
    .D(_00387_),
    .Q(\core.cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15501_ (.CLK(clk),
    .D(_00388_),
    .Q(\core.cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15502_ (.CLK(clk),
    .D(_00389_),
    .Q(\core.cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15503_ (.CLK(clk),
    .D(_00390_),
    .Q(\core.cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15504_ (.CLK(clk),
    .D(_00391_),
    .Q(\core.cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15505_ (.CLK(clk),
    .D(_00392_),
    .Q(\core.cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15506_ (.CLK(clk),
    .D(_00393_),
    .Q(\core.cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15507_ (.CLK(clk),
    .D(_00394_),
    .Q(\core.cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15508_ (.CLK(clk),
    .D(_00395_),
    .Q(\core.cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15509_ (.CLK(clk),
    .D(_00396_),
    .Q(\core.cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15510_ (.CLK(clk),
    .D(_00397_),
    .Q(\core.cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15511_ (.CLK(clk),
    .D(_00398_),
    .Q(\core.cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15512_ (.CLK(clk),
    .D(_00399_),
    .Q(\core.cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15513_ (.CLK(clk),
    .D(_00400_),
    .Q(\core.cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15514_ (.CLK(clk),
    .D(_00401_),
    .Q(\core.cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15515_ (.CLK(clk),
    .D(_00402_),
    .Q(\core.cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15516_ (.CLK(clk),
    .D(_00403_),
    .Q(\core.cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15517_ (.CLK(clk),
    .D(_00404_),
    .Q(\core.cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15518_ (.CLK(clk),
    .D(_00405_),
    .Q(\core.cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15519_ (.CLK(clk),
    .D(_00406_),
    .Q(\core.cpuregs[27][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15520_ (.CLK(clk),
    .D(_00407_),
    .Q(\core.cpuregs[27][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15521_ (.CLK(clk),
    .D(_00408_),
    .Q(\core.cpuregs[27][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15522_ (.CLK(clk),
    .D(_00409_),
    .Q(\core.cpuregs[27][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15523_ (.CLK(clk),
    .D(_00410_),
    .Q(\core.cpuregs[27][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15524_ (.CLK(clk),
    .D(_00411_),
    .Q(\core.cpuregs[27][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15525_ (.CLK(clk),
    .D(_00412_),
    .Q(\core.cpuregs[27][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15526_ (.CLK(clk),
    .D(_00413_),
    .Q(\core.cpuregs[27][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15527_ (.CLK(clk),
    .D(_00414_),
    .Q(\core.cpuregs[27][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15528_ (.CLK(clk),
    .D(_00415_),
    .Q(\core.cpuregs[27][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15529_ (.CLK(clk),
    .D(_00416_),
    .Q(\core.cpuregs[27][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15530_ (.CLK(clk),
    .D(_00417_),
    .Q(\core.cpuregs[27][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15531_ (.CLK(clk),
    .D(_00418_),
    .Q(\core.cpuregs[27][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15532_ (.CLK(clk),
    .D(_00419_),
    .Q(\core.cpuregs[27][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15533_ (.CLK(clk),
    .D(_00420_),
    .Q(\core.cpuregs[27][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15534_ (.CLK(clk),
    .D(_00421_),
    .Q(\core.cpuregs[27][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15535_ (.CLK(clk),
    .D(_00422_),
    .Q(\core.cpuregs[27][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15536_ (.CLK(clk),
    .D(_00423_),
    .Q(\core.cpuregs[27][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15537_ (.CLK(clk),
    .D(_00424_),
    .Q(\core.cpuregs[27][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15538_ (.CLK(clk),
    .D(_00425_),
    .Q(\core.cpuregs[27][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15539_ (.CLK(clk),
    .D(_00426_),
    .Q(\core.cpuregs[27][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15540_ (.CLK(clk),
    .D(_00427_),
    .Q(\core.cpuregs[27][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15541_ (.CLK(clk),
    .D(_00428_),
    .Q(\core.cpuregs[27][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15542_ (.CLK(clk),
    .D(_00429_),
    .Q(\core.cpuregs[27][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15543_ (.CLK(clk),
    .D(_00430_),
    .Q(\core.cpuregs[27][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15544_ (.CLK(clk),
    .D(_00431_),
    .Q(\core.cpuregs[27][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15545_ (.CLK(clk),
    .D(_00432_),
    .Q(\core.cpuregs[27][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15546_ (.CLK(clk),
    .D(_00433_),
    .Q(\core.cpuregs[27][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15547_ (.CLK(clk),
    .D(_00434_),
    .Q(\core.cpuregs[27][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15548_ (.CLK(clk),
    .D(_00435_),
    .Q(\core.cpuregs[27][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15549_ (.CLK(clk),
    .D(_00436_),
    .Q(\core.cpuregs[27][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15550_ (.CLK(clk),
    .D(_00437_),
    .Q(\core.cpuregs[27][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15551_ (.CLK(clk),
    .D(_00438_),
    .Q(mem_wdata[0]));
 sky130_fd_sc_hd__dfxtp_2 _15552_ (.CLK(clk),
    .D(_00439_),
    .Q(mem_wdata[1]));
 sky130_fd_sc_hd__dfxtp_2 _15553_ (.CLK(clk),
    .D(_00440_),
    .Q(mem_wdata[2]));
 sky130_fd_sc_hd__dfxtp_2 _15554_ (.CLK(clk),
    .D(_00441_),
    .Q(mem_wdata[3]));
 sky130_fd_sc_hd__dfxtp_2 _15555_ (.CLK(clk),
    .D(_00442_),
    .Q(mem_wdata[4]));
 sky130_fd_sc_hd__dfxtp_2 _15556_ (.CLK(clk),
    .D(_00443_),
    .Q(mem_wdata[5]));
 sky130_fd_sc_hd__dfxtp_2 _15557_ (.CLK(clk),
    .D(_00444_),
    .Q(mem_wdata[6]));
 sky130_fd_sc_hd__dfxtp_2 _15558_ (.CLK(clk),
    .D(_00445_),
    .Q(mem_wdata[7]));
 sky130_fd_sc_hd__dfxtp_2 _15559_ (.CLK(clk),
    .D(_00446_),
    .Q(mem_wdata[8]));
 sky130_fd_sc_hd__dfxtp_2 _15560_ (.CLK(clk),
    .D(_00447_),
    .Q(mem_wdata[9]));
 sky130_fd_sc_hd__dfxtp_2 _15561_ (.CLK(clk),
    .D(_00448_),
    .Q(mem_wdata[10]));
 sky130_fd_sc_hd__dfxtp_2 _15562_ (.CLK(clk),
    .D(_00449_),
    .Q(mem_wdata[11]));
 sky130_fd_sc_hd__dfxtp_2 _15563_ (.CLK(clk),
    .D(_00450_),
    .Q(mem_wdata[12]));
 sky130_fd_sc_hd__dfxtp_2 _15564_ (.CLK(clk),
    .D(_00451_),
    .Q(mem_wdata[13]));
 sky130_fd_sc_hd__dfxtp_2 _15565_ (.CLK(clk),
    .D(_00452_),
    .Q(mem_wdata[14]));
 sky130_fd_sc_hd__dfxtp_2 _15566_ (.CLK(clk),
    .D(_00453_),
    .Q(mem_wdata[15]));
 sky130_fd_sc_hd__dfxtp_2 _15567_ (.CLK(clk),
    .D(_00454_),
    .Q(mem_wdata[16]));
 sky130_fd_sc_hd__dfxtp_2 _15568_ (.CLK(clk),
    .D(_00455_),
    .Q(mem_wdata[17]));
 sky130_fd_sc_hd__dfxtp_2 _15569_ (.CLK(clk),
    .D(_00456_),
    .Q(mem_wdata[18]));
 sky130_fd_sc_hd__dfxtp_2 _15570_ (.CLK(clk),
    .D(_00457_),
    .Q(mem_wdata[19]));
 sky130_fd_sc_hd__dfxtp_2 _15571_ (.CLK(clk),
    .D(_00458_),
    .Q(mem_wdata[20]));
 sky130_fd_sc_hd__dfxtp_2 _15572_ (.CLK(clk),
    .D(_00459_),
    .Q(mem_wdata[21]));
 sky130_fd_sc_hd__dfxtp_2 _15573_ (.CLK(clk),
    .D(_00460_),
    .Q(mem_wdata[22]));
 sky130_fd_sc_hd__dfxtp_2 _15574_ (.CLK(clk),
    .D(_00461_),
    .Q(mem_wdata[23]));
 sky130_fd_sc_hd__dfxtp_2 _15575_ (.CLK(clk),
    .D(_00462_),
    .Q(mem_wdata[24]));
 sky130_fd_sc_hd__dfxtp_2 _15576_ (.CLK(clk),
    .D(_00463_),
    .Q(mem_wdata[25]));
 sky130_fd_sc_hd__dfxtp_2 _15577_ (.CLK(clk),
    .D(_00464_),
    .Q(mem_wdata[26]));
 sky130_fd_sc_hd__dfxtp_2 _15578_ (.CLK(clk),
    .D(_00465_),
    .Q(mem_wdata[27]));
 sky130_fd_sc_hd__dfxtp_2 _15579_ (.CLK(clk),
    .D(_00466_),
    .Q(mem_wdata[28]));
 sky130_fd_sc_hd__dfxtp_2 _15580_ (.CLK(clk),
    .D(_00467_),
    .Q(mem_wdata[29]));
 sky130_fd_sc_hd__dfxtp_2 _15581_ (.CLK(clk),
    .D(_00468_),
    .Q(mem_wdata[30]));
 sky130_fd_sc_hd__dfxtp_2 _15582_ (.CLK(clk),
    .D(_00469_),
    .Q(mem_wdata[31]));
 sky130_fd_sc_hd__dfxtp_2 _15583_ (.CLK(clk),
    .D(_00470_),
    .Q(mem_instr));
 sky130_fd_sc_hd__dfxtp_2 _15584_ (.CLK(clk),
    .D(_00471_),
    .Q(\core.cpuregs[28][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15585_ (.CLK(clk),
    .D(_00472_),
    .Q(\core.cpuregs[28][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15586_ (.CLK(clk),
    .D(_00473_),
    .Q(\core.cpuregs[28][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15587_ (.CLK(clk),
    .D(_00474_),
    .Q(\core.cpuregs[28][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15588_ (.CLK(clk),
    .D(_00475_),
    .Q(\core.cpuregs[28][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15589_ (.CLK(clk),
    .D(_00476_),
    .Q(\core.cpuregs[28][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15590_ (.CLK(clk),
    .D(_00477_),
    .Q(\core.cpuregs[28][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15591_ (.CLK(clk),
    .D(_00478_),
    .Q(\core.cpuregs[28][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15592_ (.CLK(clk),
    .D(_00479_),
    .Q(\core.cpuregs[28][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15593_ (.CLK(clk),
    .D(_00480_),
    .Q(\core.cpuregs[28][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15594_ (.CLK(clk),
    .D(_00481_),
    .Q(\core.cpuregs[28][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15595_ (.CLK(clk),
    .D(_00482_),
    .Q(\core.cpuregs[28][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15596_ (.CLK(clk),
    .D(_00483_),
    .Q(\core.cpuregs[28][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15597_ (.CLK(clk),
    .D(_00484_),
    .Q(\core.cpuregs[28][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15598_ (.CLK(clk),
    .D(_00485_),
    .Q(\core.cpuregs[28][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15599_ (.CLK(clk),
    .D(_00486_),
    .Q(\core.cpuregs[28][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15600_ (.CLK(clk),
    .D(_00487_),
    .Q(\core.cpuregs[28][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15601_ (.CLK(clk),
    .D(_00488_),
    .Q(\core.cpuregs[28][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15602_ (.CLK(clk),
    .D(_00489_),
    .Q(\core.cpuregs[28][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15603_ (.CLK(clk),
    .D(_00490_),
    .Q(\core.cpuregs[28][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15604_ (.CLK(clk),
    .D(_00491_),
    .Q(\core.cpuregs[28][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15605_ (.CLK(clk),
    .D(_00492_),
    .Q(\core.cpuregs[28][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15606_ (.CLK(clk),
    .D(_00493_),
    .Q(\core.cpuregs[28][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15607_ (.CLK(clk),
    .D(_00494_),
    .Q(\core.cpuregs[28][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15608_ (.CLK(clk),
    .D(_00495_),
    .Q(\core.cpuregs[28][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15609_ (.CLK(clk),
    .D(_00496_),
    .Q(\core.cpuregs[28][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15610_ (.CLK(clk),
    .D(_00497_),
    .Q(\core.cpuregs[28][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15611_ (.CLK(clk),
    .D(_00498_),
    .Q(\core.cpuregs[28][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15612_ (.CLK(clk),
    .D(_00499_),
    .Q(\core.cpuregs[28][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15613_ (.CLK(clk),
    .D(_00500_),
    .Q(\core.cpuregs[28][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15614_ (.CLK(clk),
    .D(_00501_),
    .Q(\core.cpuregs[28][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15615_ (.CLK(clk),
    .D(_00502_),
    .Q(\core.cpuregs[28][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15616_ (.CLK(clk),
    .D(_00503_),
    .Q(\core.is_alu_reg_reg ));
 sky130_fd_sc_hd__dfxtp_2 _15617_ (.CLK(clk),
    .D(_00504_),
    .Q(\core.is_alu_reg_imm ));
 sky130_fd_sc_hd__dfxtp_2 _15618_ (.CLK(clk),
    .D(_00505_),
    .Q(\core.instr_auipc ));
 sky130_fd_sc_hd__dfxtp_2 _15619_ (.CLK(clk),
    .D(_00506_),
    .Q(\core.instr_lui ));
 sky130_fd_sc_hd__dfxtp_2 _15620_ (.CLK(clk),
    .D(\core.alu_out[0] ),
    .Q(\core.alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15621_ (.CLK(clk),
    .D(\core.alu_out[1] ),
    .Q(\core.alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15622_ (.CLK(clk),
    .D(\core.alu_out[2] ),
    .Q(\core.alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15623_ (.CLK(clk),
    .D(\core.alu_out[3] ),
    .Q(\core.alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15624_ (.CLK(clk),
    .D(\core.alu_out[4] ),
    .Q(\core.alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15625_ (.CLK(clk),
    .D(\core.alu_out[5] ),
    .Q(\core.alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15626_ (.CLK(clk),
    .D(\core.alu_out[6] ),
    .Q(\core.alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15627_ (.CLK(clk),
    .D(\core.alu_out[7] ),
    .Q(\core.alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15628_ (.CLK(clk),
    .D(\core.alu_out[8] ),
    .Q(\core.alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15629_ (.CLK(clk),
    .D(\core.alu_out[9] ),
    .Q(\core.alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15630_ (.CLK(clk),
    .D(\core.alu_out[10] ),
    .Q(\core.alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15631_ (.CLK(clk),
    .D(\core.alu_out[11] ),
    .Q(\core.alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15632_ (.CLK(clk),
    .D(\core.alu_out[12] ),
    .Q(\core.alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15633_ (.CLK(clk),
    .D(\core.alu_out[13] ),
    .Q(\core.alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15634_ (.CLK(clk),
    .D(\core.alu_out[14] ),
    .Q(\core.alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15635_ (.CLK(clk),
    .D(\core.alu_out[15] ),
    .Q(\core.alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15636_ (.CLK(clk),
    .D(\core.alu_out[16] ),
    .Q(\core.alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15637_ (.CLK(clk),
    .D(\core.alu_out[17] ),
    .Q(\core.alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15638_ (.CLK(clk),
    .D(\core.alu_out[18] ),
    .Q(\core.alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15639_ (.CLK(clk),
    .D(\core.alu_out[19] ),
    .Q(\core.alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15640_ (.CLK(clk),
    .D(\core.alu_out[20] ),
    .Q(\core.alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15641_ (.CLK(clk),
    .D(\core.alu_out[21] ),
    .Q(\core.alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15642_ (.CLK(clk),
    .D(\core.alu_out[22] ),
    .Q(\core.alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15643_ (.CLK(clk),
    .D(\core.alu_out[23] ),
    .Q(\core.alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15644_ (.CLK(clk),
    .D(\core.alu_out[24] ),
    .Q(\core.alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15645_ (.CLK(clk),
    .D(\core.alu_out[25] ),
    .Q(\core.alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15646_ (.CLK(clk),
    .D(\core.alu_out[26] ),
    .Q(\core.alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15647_ (.CLK(clk),
    .D(\core.alu_out[27] ),
    .Q(\core.alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15648_ (.CLK(clk),
    .D(\core.alu_out[28] ),
    .Q(\core.alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15649_ (.CLK(clk),
    .D(\core.alu_out[29] ),
    .Q(\core.alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15650_ (.CLK(clk),
    .D(\core.alu_out[30] ),
    .Q(\core.alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15651_ (.CLK(clk),
    .D(\core.alu_out[31] ),
    .Q(\core.alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15652_ (.CLK(clk),
    .D(_00507_),
    .Q(\core.latched_is_lb ));
 sky130_fd_sc_hd__dfxtp_2 _15653_ (.CLK(clk),
    .D(_00508_),
    .Q(\core.latched_is_lh ));
 sky130_fd_sc_hd__dfxtp_2 _15654_ (.CLK(clk),
    .D(_00509_),
    .Q(\core.decoder_pseudo_trigger ));
 sky130_fd_sc_hd__dfxtp_2 _15655_ (.CLK(clk),
    .D(_00510_),
    .Q(\core.latched_branch ));
 sky130_fd_sc_hd__dfxtp_2 _15656_ (.CLK(clk),
    .D(_00511_),
    .Q(\core.latched_stalu ));
 sky130_fd_sc_hd__dfxtp_2 _15657_ (.CLK(clk),
    .D(_00512_),
    .Q(trap));
 sky130_fd_sc_hd__dfxtp_2 _15658_ (.CLK(clk),
    .D(_00513_),
    .Q(\core.instr_bne ));
 sky130_fd_sc_hd__dfxtp_2 _15659_ (.CLK(clk),
    .D(_00514_),
    .Q(\core.cpuregs[21][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15660_ (.CLK(clk),
    .D(_00515_),
    .Q(\core.cpuregs[21][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15661_ (.CLK(clk),
    .D(_00516_),
    .Q(\core.cpuregs[21][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15662_ (.CLK(clk),
    .D(_00517_),
    .Q(\core.cpuregs[21][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15663_ (.CLK(clk),
    .D(_00518_),
    .Q(\core.cpuregs[21][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15664_ (.CLK(clk),
    .D(_00519_),
    .Q(\core.cpuregs[21][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15665_ (.CLK(clk),
    .D(_00520_),
    .Q(\core.cpuregs[21][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15666_ (.CLK(clk),
    .D(_00521_),
    .Q(\core.cpuregs[21][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15667_ (.CLK(clk),
    .D(_00522_),
    .Q(\core.cpuregs[21][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15668_ (.CLK(clk),
    .D(_00523_),
    .Q(\core.cpuregs[21][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15669_ (.CLK(clk),
    .D(_00524_),
    .Q(\core.cpuregs[21][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15670_ (.CLK(clk),
    .D(_00525_),
    .Q(\core.cpuregs[21][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15671_ (.CLK(clk),
    .D(_00526_),
    .Q(\core.cpuregs[21][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15672_ (.CLK(clk),
    .D(_00527_),
    .Q(\core.cpuregs[21][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15673_ (.CLK(clk),
    .D(_00528_),
    .Q(\core.cpuregs[21][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15674_ (.CLK(clk),
    .D(_00529_),
    .Q(\core.cpuregs[21][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15675_ (.CLK(clk),
    .D(_00530_),
    .Q(\core.cpuregs[21][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15676_ (.CLK(clk),
    .D(_00531_),
    .Q(\core.cpuregs[21][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15677_ (.CLK(clk),
    .D(_00532_),
    .Q(\core.cpuregs[21][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15678_ (.CLK(clk),
    .D(_00533_),
    .Q(\core.cpuregs[21][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15679_ (.CLK(clk),
    .D(_00534_),
    .Q(\core.cpuregs[21][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15680_ (.CLK(clk),
    .D(_00535_),
    .Q(\core.cpuregs[21][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15681_ (.CLK(clk),
    .D(_00536_),
    .Q(\core.cpuregs[21][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15682_ (.CLK(clk),
    .D(_00537_),
    .Q(\core.cpuregs[21][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15683_ (.CLK(clk),
    .D(_00538_),
    .Q(\core.cpuregs[21][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15684_ (.CLK(clk),
    .D(_00539_),
    .Q(\core.cpuregs[21][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15685_ (.CLK(clk),
    .D(_00540_),
    .Q(\core.cpuregs[21][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15686_ (.CLK(clk),
    .D(_00541_),
    .Q(\core.cpuregs[21][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15687_ (.CLK(clk),
    .D(_00542_),
    .Q(\core.cpuregs[21][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15688_ (.CLK(clk),
    .D(_00543_),
    .Q(\core.cpuregs[21][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15689_ (.CLK(clk),
    .D(_00544_),
    .Q(\core.cpuregs[21][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15690_ (.CLK(clk),
    .D(_00545_),
    .Q(\core.cpuregs[21][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15691_ (.CLK(clk),
    .D(_00546_),
    .Q(\core.instr_jal ));
 sky130_fd_sc_hd__dfxtp_2 _15692_ (.CLK(clk),
    .D(_00547_),
    .Q(\core.instr_beq ));
 sky130_fd_sc_hd__dfxtp_2 _15693_ (.CLK(clk),
    .D(_00548_),
    .Q(\core.cpuregs[26][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15694_ (.CLK(clk),
    .D(_00549_),
    .Q(\core.cpuregs[26][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15695_ (.CLK(clk),
    .D(_00550_),
    .Q(\core.cpuregs[26][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15696_ (.CLK(clk),
    .D(_00551_),
    .Q(\core.cpuregs[26][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15697_ (.CLK(clk),
    .D(_00552_),
    .Q(\core.cpuregs[26][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15698_ (.CLK(clk),
    .D(_00553_),
    .Q(\core.cpuregs[26][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15699_ (.CLK(clk),
    .D(_00554_),
    .Q(\core.cpuregs[26][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15700_ (.CLK(clk),
    .D(_00555_),
    .Q(\core.cpuregs[26][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15701_ (.CLK(clk),
    .D(_00556_),
    .Q(\core.cpuregs[26][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15702_ (.CLK(clk),
    .D(_00557_),
    .Q(\core.cpuregs[26][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15703_ (.CLK(clk),
    .D(_00558_),
    .Q(\core.cpuregs[26][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15704_ (.CLK(clk),
    .D(_00559_),
    .Q(\core.cpuregs[26][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15705_ (.CLK(clk),
    .D(_00560_),
    .Q(\core.cpuregs[26][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15706_ (.CLK(clk),
    .D(_00561_),
    .Q(\core.cpuregs[26][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15707_ (.CLK(clk),
    .D(_00562_),
    .Q(\core.cpuregs[26][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15708_ (.CLK(clk),
    .D(_00563_),
    .Q(\core.cpuregs[26][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15709_ (.CLK(clk),
    .D(_00564_),
    .Q(\core.cpuregs[26][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15710_ (.CLK(clk),
    .D(_00565_),
    .Q(\core.cpuregs[26][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15711_ (.CLK(clk),
    .D(_00566_),
    .Q(\core.cpuregs[26][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15712_ (.CLK(clk),
    .D(_00567_),
    .Q(\core.cpuregs[26][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15713_ (.CLK(clk),
    .D(_00568_),
    .Q(\core.cpuregs[26][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15714_ (.CLK(clk),
    .D(_00569_),
    .Q(\core.cpuregs[26][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15715_ (.CLK(clk),
    .D(_00570_),
    .Q(\core.cpuregs[26][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15716_ (.CLK(clk),
    .D(_00571_),
    .Q(\core.cpuregs[26][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15717_ (.CLK(clk),
    .D(_00572_),
    .Q(\core.cpuregs[26][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15718_ (.CLK(clk),
    .D(_00573_),
    .Q(\core.cpuregs[26][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15719_ (.CLK(clk),
    .D(_00574_),
    .Q(\core.cpuregs[26][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15720_ (.CLK(clk),
    .D(_00575_),
    .Q(\core.cpuregs[26][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15721_ (.CLK(clk),
    .D(_00576_),
    .Q(\core.cpuregs[26][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15722_ (.CLK(clk),
    .D(_00577_),
    .Q(\core.cpuregs[26][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15723_ (.CLK(clk),
    .D(_00578_),
    .Q(\core.cpuregs[26][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15724_ (.CLK(clk),
    .D(_00579_),
    .Q(\core.cpuregs[26][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15725_ (.CLK(clk),
    .D(_00580_),
    .Q(\core.instr_sh ));
 sky130_fd_sc_hd__dfxtp_2 _15726_ (.CLK(clk),
    .D(_00581_),
    .Q(\core.instr_slti ));
 sky130_fd_sc_hd__dfxtp_2 _15727_ (.CLK(clk),
    .D(_00582_),
    .Q(\core.instr_sltiu ));
 sky130_fd_sc_hd__dfxtp_2 _15728_ (.CLK(clk),
    .D(_00583_),
    .Q(\core.instr_ori ));
 sky130_fd_sc_hd__dfxtp_2 _15729_ (.CLK(clk),
    .D(_00584_),
    .Q(\core.latched_store ));
 sky130_fd_sc_hd__dfxtp_2 _15730_ (.CLK(clk),
    .D(_00585_),
    .Q(\core.instr_srli ));
 sky130_fd_sc_hd__dfxtp_2 _15731_ (.CLK(clk),
    .D(_00586_),
    .Q(\core.instr_add ));
 sky130_fd_sc_hd__dfxtp_2 _15732_ (.CLK(clk),
    .D(_00587_),
    .Q(\core.instr_sll ));
 sky130_fd_sc_hd__dfxtp_2 _15733_ (.CLK(clk),
    .D(_00588_),
    .Q(\core.instr_xor ));
 sky130_fd_sc_hd__dfxtp_2 _15734_ (.CLK(clk),
    .D(_00589_),
    .Q(\core.instr_sra ));
 sky130_fd_sc_hd__dfxtp_2 _15735_ (.CLK(clk),
    .D(_00590_),
    .Q(\core.is_compare ));
 sky130_fd_sc_hd__dfxtp_2 _15736_ (.CLK(clk),
    .D(_00591_),
    .Q(\core.latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15737_ (.CLK(clk),
    .D(_00592_),
    .Q(\core.latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15738_ (.CLK(clk),
    .D(_00593_),
    .Q(\core.latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15739_ (.CLK(clk),
    .D(_00594_),
    .Q(\core.latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15740_ (.CLK(clk),
    .D(_00595_),
    .Q(\core.latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15741_ (.CLK(clk),
    .D(_00596_),
    .Q(mem_wstrb[0]));
 sky130_fd_sc_hd__dfxtp_2 _15742_ (.CLK(clk),
    .D(_00597_),
    .Q(mem_wstrb[1]));
 sky130_fd_sc_hd__dfxtp_2 _15743_ (.CLK(clk),
    .D(_00598_),
    .Q(mem_wstrb[2]));
 sky130_fd_sc_hd__dfxtp_2 _15744_ (.CLK(clk),
    .D(_00599_),
    .Q(mem_wstrb[3]));
 sky130_fd_sc_hd__dfxtp_2 _15745_ (.CLK(clk),
    .D(_00600_),
    .Q(\core.instr_rdcycleh ));
 sky130_fd_sc_hd__dfxtp_2 _15746_ (.CLK(clk),
    .D(_00601_),
    .Q(mem_valid));
 sky130_fd_sc_hd__dfxtp_2 _15747_ (.CLK(clk),
    .D(_00602_),
    .Q(\core.instr_fence ));
 sky130_fd_sc_hd__dfxtp_2 _15748_ (.CLK(clk),
    .D(_00603_),
    .Q(\core.mem_do_wdata ));
 sky130_fd_sc_hd__dfxtp_2 _15749_ (.CLK(clk),
    .D(_00030_),
    .Q(\core.decoder_trigger ));
 sky130_fd_sc_hd__dfxtp_2 _15750_ (.CLK(clk),
    .D(_00604_),
    .Q(\core.mem_la_wdata[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15751_ (.CLK(clk),
    .D(_00605_),
    .Q(\core.mem_la_wdata[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15752_ (.CLK(clk),
    .D(_00606_),
    .Q(\core.mem_la_wdata[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15753_ (.CLK(clk),
    .D(_00607_),
    .Q(\core.mem_la_wdata[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15754_ (.CLK(clk),
    .D(_00608_),
    .Q(\core.mem_la_wdata[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15755_ (.CLK(clk),
    .D(_00609_),
    .Q(\core.mem_la_wdata[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15756_ (.CLK(clk),
    .D(_00610_),
    .Q(\core.mem_la_wdata[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15757_ (.CLK(clk),
    .D(_00611_),
    .Q(\core.mem_la_wdata[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15758_ (.CLK(clk),
    .D(_00612_),
    .Q(\core.pcpi_rs2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15759_ (.CLK(clk),
    .D(_00613_),
    .Q(\core.pcpi_rs2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15760_ (.CLK(clk),
    .D(_00614_),
    .Q(\core.pcpi_rs2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15761_ (.CLK(clk),
    .D(_00615_),
    .Q(\core.pcpi_rs2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15762_ (.CLK(clk),
    .D(_00616_),
    .Q(\core.pcpi_rs2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15763_ (.CLK(clk),
    .D(_00617_),
    .Q(\core.pcpi_rs2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15764_ (.CLK(clk),
    .D(_00618_),
    .Q(\core.pcpi_rs2[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15765_ (.CLK(clk),
    .D(_00619_),
    .Q(\core.pcpi_rs2[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15766_ (.CLK(clk),
    .D(_00620_),
    .Q(\core.pcpi_rs2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15767_ (.CLK(clk),
    .D(_00621_),
    .Q(\core.pcpi_rs2[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15768_ (.CLK(clk),
    .D(_00622_),
    .Q(\core.pcpi_rs2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15769_ (.CLK(clk),
    .D(_00623_),
    .Q(\core.pcpi_rs2[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15770_ (.CLK(clk),
    .D(_00624_),
    .Q(\core.pcpi_rs2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15771_ (.CLK(clk),
    .D(_00625_),
    .Q(\core.pcpi_rs2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15772_ (.CLK(clk),
    .D(_00626_),
    .Q(\core.pcpi_rs2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15773_ (.CLK(clk),
    .D(_00627_),
    .Q(\core.pcpi_rs2[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15774_ (.CLK(clk),
    .D(_00628_),
    .Q(\core.pcpi_rs2[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15775_ (.CLK(clk),
    .D(_00629_),
    .Q(\core.pcpi_rs2[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15776_ (.CLK(clk),
    .D(_00630_),
    .Q(\core.pcpi_rs2[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15777_ (.CLK(clk),
    .D(_00631_),
    .Q(\core.pcpi_rs2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15778_ (.CLK(clk),
    .D(_00632_),
    .Q(\core.pcpi_rs2[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15779_ (.CLK(clk),
    .D(_00633_),
    .Q(\core.pcpi_rs2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15780_ (.CLK(clk),
    .D(_00634_),
    .Q(\core.pcpi_rs2[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15781_ (.CLK(clk),
    .D(_00635_),
    .Q(\core.pcpi_rs2[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15782_ (.CLK(clk),
    .D(_00636_),
    .Q(\core.instr_bge ));
 sky130_fd_sc_hd__dfxtp_2 _15783_ (.CLK(clk),
    .D(_00637_),
    .Q(\core.instr_bltu ));
 sky130_fd_sc_hd__dfxtp_2 _15784_ (.CLK(clk),
    .D(_00638_),
    .Q(\core.instr_jalr ));
 sky130_fd_sc_hd__dfxtp_2 _15785_ (.CLK(clk),
    .D(_00639_),
    .Q(\core.instr_lb ));
 sky130_fd_sc_hd__dfxtp_2 _15786_ (.CLK(clk),
    .D(_00640_),
    .Q(\core.cpuregs[20][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15787_ (.CLK(clk),
    .D(_00641_),
    .Q(\core.cpuregs[20][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15788_ (.CLK(clk),
    .D(_00642_),
    .Q(\core.cpuregs[20][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15789_ (.CLK(clk),
    .D(_00643_),
    .Q(\core.cpuregs[20][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15790_ (.CLK(clk),
    .D(_00644_),
    .Q(\core.cpuregs[20][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15791_ (.CLK(clk),
    .D(_00645_),
    .Q(\core.cpuregs[20][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15792_ (.CLK(clk),
    .D(_00646_),
    .Q(\core.cpuregs[20][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15793_ (.CLK(clk),
    .D(_00647_),
    .Q(\core.cpuregs[20][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15794_ (.CLK(clk),
    .D(_00648_),
    .Q(\core.cpuregs[20][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15795_ (.CLK(clk),
    .D(_00649_),
    .Q(\core.cpuregs[20][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15796_ (.CLK(clk),
    .D(_00650_),
    .Q(\core.cpuregs[20][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15797_ (.CLK(clk),
    .D(_00651_),
    .Q(\core.cpuregs[20][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15798_ (.CLK(clk),
    .D(_00652_),
    .Q(\core.cpuregs[20][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15799_ (.CLK(clk),
    .D(_00653_),
    .Q(\core.cpuregs[20][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15800_ (.CLK(clk),
    .D(_00654_),
    .Q(\core.cpuregs[20][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15801_ (.CLK(clk),
    .D(_00655_),
    .Q(\core.cpuregs[20][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15802_ (.CLK(clk),
    .D(_00656_),
    .Q(\core.cpuregs[20][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15803_ (.CLK(clk),
    .D(_00657_),
    .Q(\core.cpuregs[20][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15804_ (.CLK(clk),
    .D(_00658_),
    .Q(\core.cpuregs[20][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15805_ (.CLK(clk),
    .D(_00659_),
    .Q(\core.cpuregs[20][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15806_ (.CLK(clk),
    .D(_00660_),
    .Q(\core.cpuregs[20][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15807_ (.CLK(clk),
    .D(_00661_),
    .Q(\core.cpuregs[20][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15808_ (.CLK(clk),
    .D(_00662_),
    .Q(\core.cpuregs[20][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15809_ (.CLK(clk),
    .D(_00663_),
    .Q(\core.cpuregs[20][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15810_ (.CLK(clk),
    .D(_00664_),
    .Q(\core.cpuregs[20][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15811_ (.CLK(clk),
    .D(_00665_),
    .Q(\core.cpuregs[20][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15812_ (.CLK(clk),
    .D(_00666_),
    .Q(\core.cpuregs[20][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15813_ (.CLK(clk),
    .D(_00667_),
    .Q(\core.cpuregs[20][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15814_ (.CLK(clk),
    .D(_00668_),
    .Q(\core.cpuregs[20][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15815_ (.CLK(clk),
    .D(_00669_),
    .Q(\core.cpuregs[20][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15816_ (.CLK(clk),
    .D(_00670_),
    .Q(\core.cpuregs[20][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15817_ (.CLK(clk),
    .D(_00671_),
    .Q(\core.cpuregs[20][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15818_ (.CLK(clk),
    .D(_00672_),
    .Q(\core.cpuregs[25][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15819_ (.CLK(clk),
    .D(_00673_),
    .Q(\core.cpuregs[25][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15820_ (.CLK(clk),
    .D(_00674_),
    .Q(\core.cpuregs[25][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15821_ (.CLK(clk),
    .D(_00675_),
    .Q(\core.cpuregs[25][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15822_ (.CLK(clk),
    .D(_00676_),
    .Q(\core.cpuregs[25][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15823_ (.CLK(clk),
    .D(_00677_),
    .Q(\core.cpuregs[25][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15824_ (.CLK(clk),
    .D(_00678_),
    .Q(\core.cpuregs[25][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15825_ (.CLK(clk),
    .D(_00679_),
    .Q(\core.cpuregs[25][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15826_ (.CLK(clk),
    .D(_00680_),
    .Q(\core.cpuregs[25][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15827_ (.CLK(clk),
    .D(_00681_),
    .Q(\core.cpuregs[25][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15828_ (.CLK(clk),
    .D(_00682_),
    .Q(\core.cpuregs[25][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15829_ (.CLK(clk),
    .D(_00683_),
    .Q(\core.cpuregs[25][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15830_ (.CLK(clk),
    .D(_00684_),
    .Q(\core.cpuregs[25][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15831_ (.CLK(clk),
    .D(_00685_),
    .Q(\core.cpuregs[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15832_ (.CLK(clk),
    .D(_00686_),
    .Q(\core.cpuregs[25][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15833_ (.CLK(clk),
    .D(_00687_),
    .Q(\core.cpuregs[25][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15834_ (.CLK(clk),
    .D(_00688_),
    .Q(\core.cpuregs[25][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15835_ (.CLK(clk),
    .D(_00689_),
    .Q(\core.cpuregs[25][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15836_ (.CLK(clk),
    .D(_00690_),
    .Q(\core.cpuregs[25][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15837_ (.CLK(clk),
    .D(_00691_),
    .Q(\core.cpuregs[25][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15838_ (.CLK(clk),
    .D(_00692_),
    .Q(\core.cpuregs[25][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15839_ (.CLK(clk),
    .D(_00693_),
    .Q(\core.cpuregs[25][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15840_ (.CLK(clk),
    .D(_00694_),
    .Q(\core.cpuregs[25][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15841_ (.CLK(clk),
    .D(_00695_),
    .Q(\core.cpuregs[25][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15842_ (.CLK(clk),
    .D(_00696_),
    .Q(\core.cpuregs[25][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15843_ (.CLK(clk),
    .D(_00697_),
    .Q(\core.cpuregs[25][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15844_ (.CLK(clk),
    .D(_00698_),
    .Q(\core.cpuregs[25][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15845_ (.CLK(clk),
    .D(_00699_),
    .Q(\core.cpuregs[25][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15846_ (.CLK(clk),
    .D(_00700_),
    .Q(\core.cpuregs[25][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15847_ (.CLK(clk),
    .D(_00701_),
    .Q(\core.cpuregs[25][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15848_ (.CLK(clk),
    .D(_00702_),
    .Q(\core.cpuregs[25][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15849_ (.CLK(clk),
    .D(_00703_),
    .Q(\core.cpuregs[25][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15850_ (.CLK(clk),
    .D(_00704_),
    .Q(\core.cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15851_ (.CLK(clk),
    .D(_00705_),
    .Q(\core.cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15852_ (.CLK(clk),
    .D(_00706_),
    .Q(\core.cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15853_ (.CLK(clk),
    .D(_00707_),
    .Q(\core.cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15854_ (.CLK(clk),
    .D(_00708_),
    .Q(\core.cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15855_ (.CLK(clk),
    .D(_00709_),
    .Q(\core.cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15856_ (.CLK(clk),
    .D(_00710_),
    .Q(\core.cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15857_ (.CLK(clk),
    .D(_00711_),
    .Q(\core.cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15858_ (.CLK(clk),
    .D(_00712_),
    .Q(\core.cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15859_ (.CLK(clk),
    .D(_00713_),
    .Q(\core.cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15860_ (.CLK(clk),
    .D(_00714_),
    .Q(\core.cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15861_ (.CLK(clk),
    .D(_00715_),
    .Q(\core.cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15862_ (.CLK(clk),
    .D(_00716_),
    .Q(\core.cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15863_ (.CLK(clk),
    .D(_00717_),
    .Q(\core.cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15864_ (.CLK(clk),
    .D(_00718_),
    .Q(\core.cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15865_ (.CLK(clk),
    .D(_00719_),
    .Q(\core.cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15866_ (.CLK(clk),
    .D(_00720_),
    .Q(\core.cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15867_ (.CLK(clk),
    .D(_00721_),
    .Q(\core.cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15868_ (.CLK(clk),
    .D(_00722_),
    .Q(\core.cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15869_ (.CLK(clk),
    .D(_00723_),
    .Q(\core.cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15870_ (.CLK(clk),
    .D(_00724_),
    .Q(\core.cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15871_ (.CLK(clk),
    .D(_00725_),
    .Q(\core.cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15872_ (.CLK(clk),
    .D(_00726_),
    .Q(\core.cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15873_ (.CLK(clk),
    .D(_00727_),
    .Q(\core.cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15874_ (.CLK(clk),
    .D(_00728_),
    .Q(\core.cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15875_ (.CLK(clk),
    .D(_00729_),
    .Q(\core.cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15876_ (.CLK(clk),
    .D(_00730_),
    .Q(\core.cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15877_ (.CLK(clk),
    .D(_00731_),
    .Q(\core.cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15878_ (.CLK(clk),
    .D(_00732_),
    .Q(\core.cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15879_ (.CLK(clk),
    .D(_00733_),
    .Q(\core.cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15880_ (.CLK(clk),
    .D(_00734_),
    .Q(\core.cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15881_ (.CLK(clk),
    .D(_00735_),
    .Q(\core.cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15882_ (.CLK(clk),
    .D(_00736_),
    .Q(\core.decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15883_ (.CLK(clk),
    .D(_00737_),
    .Q(\core.decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15884_ (.CLK(clk),
    .D(_00738_),
    .Q(\core.decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15885_ (.CLK(clk),
    .D(_00739_),
    .Q(\core.decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15886_ (.CLK(clk),
    .D(_00740_),
    .Q(\core.decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15887_ (.CLK(clk),
    .D(_00741_),
    .Q(\core.decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_2 _15888_ (.CLK(clk),
    .D(_00031_),
    .Q(\core.is_lui_auipc_jal ));
 sky130_fd_sc_hd__dfxtp_2 _15889_ (.CLK(clk),
    .D(_00742_),
    .Q(\core.decoded_imm_j[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15890_ (.CLK(clk),
    .D(_00743_),
    .Q(\core.decoded_imm_j[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15891_ (.CLK(clk),
    .D(_00744_),
    .Q(\core.decoded_imm_j[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15892_ (.CLK(clk),
    .D(_00745_),
    .Q(\core.decoded_imm_j[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15893_ (.CLK(clk),
    .D(_00746_),
    .Q(\core.decoded_imm_j[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15894_ (.CLK(clk),
    .D(_00747_),
    .Q(\core.decoded_imm_j[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15895_ (.CLK(clk),
    .D(_00748_),
    .Q(\core.decoded_imm_j[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15896_ (.CLK(clk),
    .D(_00749_),
    .Q(\core.decoded_imm_j[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15897_ (.CLK(clk),
    .D(_00750_),
    .Q(\core.decoded_imm_j[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15898_ (.CLK(clk),
    .D(_00751_),
    .Q(\core.decoded_imm_j[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15899_ (.CLK(clk),
    .D(_00752_),
    .Q(\core.decoded_imm_j[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15900_ (.CLK(clk),
    .D(_00753_),
    .Q(\core.decoded_imm_j[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15901_ (.CLK(clk),
    .D(_00754_),
    .Q(\core.decoded_imm_j[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15902_ (.CLK(clk),
    .D(_00755_),
    .Q(\core.decoded_imm_j[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15903_ (.CLK(clk),
    .D(_00756_),
    .Q(\core.decoded_imm_j[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15904_ (.CLK(clk),
    .D(_00757_),
    .Q(\core.decoded_imm_j[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15905_ (.CLK(clk),
    .D(_00758_),
    .Q(\core.decoded_imm_j[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15906_ (.CLK(clk),
    .D(_00759_),
    .Q(\core.decoded_imm_j[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15907_ (.CLK(clk),
    .D(_00760_),
    .Q(\core.decoded_imm_j[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15908_ (.CLK(clk),
    .D(_00761_),
    .Q(\core.decoded_imm_j[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15909_ (.CLK(clk),
    .D(_00762_),
    .Q(\core.is_lb_lh_lw_lbu_lhu ));
 sky130_fd_sc_hd__dfxtp_2 _15910_ (.CLK(clk),
    .D(_00763_),
    .Q(\core.is_slli_srli_srai ));
 sky130_fd_sc_hd__dfxtp_2 _15911_ (.CLK(clk),
    .D(_00764_),
    .Q(\core.is_jalr_addi_slti_sltiu_xori_ori_andi ));
 sky130_fd_sc_hd__dfxtp_2 _15912_ (.CLK(clk),
    .D(_00765_),
    .Q(\core.is_sb_sh_sw ));
 sky130_fd_sc_hd__dfxtp_2 _15913_ (.CLK(clk),
    .D(_00766_),
    .Q(\core.is_sll_srl_sra ));
 sky130_fd_sc_hd__dfxtp_2 _15914_ (.CLK(clk),
    .D(_00032_),
    .Q(\core.is_slti_blt_slt ));
 sky130_fd_sc_hd__dfxtp_2 _15915_ (.CLK(clk),
    .D(_00033_),
    .Q(\core.is_sltiu_bltu_sltu ));
 sky130_fd_sc_hd__dfxtp_2 _15916_ (.CLK(clk),
    .D(_00767_),
    .Q(\core.is_beq_bne_blt_bge_bltu_bgeu ));
 sky130_fd_sc_hd__dfxtp_2 _15917_ (.CLK(clk),
    .D(_00768_),
    .Q(\core.decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_2 _15918_ (.CLK(clk),
    .D(_00769_),
    .Q(\core.decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15919_ (.CLK(clk),
    .D(_00770_),
    .Q(\core.decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_2 _15920_ (.CLK(clk),
    .D(_00771_),
    .Q(\core.decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15921_ (.CLK(clk),
    .D(_00772_),
    .Q(\core.decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15922_ (.CLK(clk),
    .D(_00773_),
    .Q(\core.decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15923_ (.CLK(clk),
    .D(_00774_),
    .Q(\core.decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15924_ (.CLK(clk),
    .D(_00775_),
    .Q(\core.decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15925_ (.CLK(clk),
    .D(_00776_),
    .Q(\core.decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15926_ (.CLK(clk),
    .D(_00777_),
    .Q(\core.decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15927_ (.CLK(clk),
    .D(_00778_),
    .Q(\core.decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15928_ (.CLK(clk),
    .D(_00779_),
    .Q(\core.decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15929_ (.CLK(clk),
    .D(_00780_),
    .Q(\core.decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15930_ (.CLK(clk),
    .D(_00781_),
    .Q(\core.decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15931_ (.CLK(clk),
    .D(_00782_),
    .Q(\core.decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15932_ (.CLK(clk),
    .D(_00783_),
    .Q(\core.decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15933_ (.CLK(clk),
    .D(_00784_),
    .Q(\core.decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15934_ (.CLK(clk),
    .D(_00785_),
    .Q(\core.decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15935_ (.CLK(clk),
    .D(_00786_),
    .Q(\core.decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 _15936_ (.CLK(clk),
    .D(_00787_),
    .Q(\core.decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _15937_ (.CLK(clk),
    .D(_00788_),
    .Q(\core.decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_2 _15938_ (.CLK(clk),
    .D(_00789_),
    .Q(\core.decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_2 _15939_ (.CLK(clk),
    .D(_00790_),
    .Q(\core.decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 _15940_ (.CLK(clk),
    .D(_00791_),
    .Q(\core.decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_2 _15941_ (.CLK(clk),
    .D(_00792_),
    .Q(\core.decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 _15942_ (.CLK(clk),
    .D(_00793_),
    .Q(\core.decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15943_ (.CLK(clk),
    .D(_00794_),
    .Q(\core.decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_2 _15944_ (.CLK(clk),
    .D(_00795_),
    .Q(\core.decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_2 _15945_ (.CLK(clk),
    .D(_00796_),
    .Q(\core.decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _15946_ (.CLK(clk),
    .D(_00797_),
    .Q(\core.decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15947_ (.CLK(clk),
    .D(_00798_),
    .Q(\core.decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_2 _15948_ (.CLK(clk),
    .D(_00799_),
    .Q(\core.cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15949_ (.CLK(clk),
    .D(_00800_),
    .Q(\core.cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15950_ (.CLK(clk),
    .D(_00801_),
    .Q(\core.cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15951_ (.CLK(clk),
    .D(_00802_),
    .Q(\core.cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15952_ (.CLK(clk),
    .D(_00803_),
    .Q(\core.cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15953_ (.CLK(clk),
    .D(_00804_),
    .Q(\core.cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15954_ (.CLK(clk),
    .D(_00805_),
    .Q(\core.cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15955_ (.CLK(clk),
    .D(_00806_),
    .Q(\core.cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15956_ (.CLK(clk),
    .D(_00807_),
    .Q(\core.cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15957_ (.CLK(clk),
    .D(_00808_),
    .Q(\core.cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15958_ (.CLK(clk),
    .D(_00809_),
    .Q(\core.cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15959_ (.CLK(clk),
    .D(_00810_),
    .Q(\core.cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15960_ (.CLK(clk),
    .D(_00811_),
    .Q(\core.cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15961_ (.CLK(clk),
    .D(_00812_),
    .Q(\core.cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15962_ (.CLK(clk),
    .D(_00813_),
    .Q(\core.cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15963_ (.CLK(clk),
    .D(_00814_),
    .Q(\core.cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15964_ (.CLK(clk),
    .D(_00815_),
    .Q(\core.cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15965_ (.CLK(clk),
    .D(_00816_),
    .Q(\core.cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15966_ (.CLK(clk),
    .D(_00817_),
    .Q(\core.cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15967_ (.CLK(clk),
    .D(_00818_),
    .Q(\core.cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _15968_ (.CLK(clk),
    .D(_00819_),
    .Q(\core.cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _15969_ (.CLK(clk),
    .D(_00820_),
    .Q(\core.cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 _15970_ (.CLK(clk),
    .D(_00821_),
    .Q(\core.cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 _15971_ (.CLK(clk),
    .D(_00822_),
    .Q(\core.cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 _15972_ (.CLK(clk),
    .D(_00823_),
    .Q(\core.cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _15973_ (.CLK(clk),
    .D(_00824_),
    .Q(\core.cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _15974_ (.CLK(clk),
    .D(_00825_),
    .Q(\core.cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _15975_ (.CLK(clk),
    .D(_00826_),
    .Q(\core.cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 _15976_ (.CLK(clk),
    .D(_00827_),
    .Q(\core.cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 _15977_ (.CLK(clk),
    .D(_00828_),
    .Q(\core.cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _15978_ (.CLK(clk),
    .D(_00829_),
    .Q(\core.cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 _15979_ (.CLK(clk),
    .D(_00830_),
    .Q(\core.cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15980_ (.CLK(clk),
    .D(_00831_),
    .Q(\core.cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _15981_ (.CLK(clk),
    .D(_00832_),
    .Q(\core.cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _15982_ (.CLK(clk),
    .D(_00833_),
    .Q(\core.cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _15983_ (.CLK(clk),
    .D(_00834_),
    .Q(\core.cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _15984_ (.CLK(clk),
    .D(_00835_),
    .Q(\core.cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _15985_ (.CLK(clk),
    .D(_00836_),
    .Q(\core.cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _15986_ (.CLK(clk),
    .D(_00837_),
    .Q(\core.cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _15987_ (.CLK(clk),
    .D(_00838_),
    .Q(\core.cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _15988_ (.CLK(clk),
    .D(_00839_),
    .Q(\core.cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 _15989_ (.CLK(clk),
    .D(_00840_),
    .Q(\core.cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 _15990_ (.CLK(clk),
    .D(_00841_),
    .Q(\core.cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _15991_ (.CLK(clk),
    .D(_00842_),
    .Q(\core.cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _15992_ (.CLK(clk),
    .D(_00843_),
    .Q(\core.cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _15993_ (.CLK(clk),
    .D(_00844_),
    .Q(\core.cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 _15994_ (.CLK(clk),
    .D(_00845_),
    .Q(\core.cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 _15995_ (.CLK(clk),
    .D(_00846_),
    .Q(\core.cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _15996_ (.CLK(clk),
    .D(_00847_),
    .Q(\core.cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 _15997_ (.CLK(clk),
    .D(_00848_),
    .Q(\core.cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 _15998_ (.CLK(clk),
    .D(_00849_),
    .Q(\core.cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 _15999_ (.CLK(clk),
    .D(_00850_),
    .Q(\core.cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16000_ (.CLK(clk),
    .D(_00851_),
    .Q(\core.cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16001_ (.CLK(clk),
    .D(_00852_),
    .Q(\core.cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16002_ (.CLK(clk),
    .D(_00853_),
    .Q(\core.cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16003_ (.CLK(clk),
    .D(_00854_),
    .Q(\core.cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16004_ (.CLK(clk),
    .D(_00855_),
    .Q(\core.cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16005_ (.CLK(clk),
    .D(_00856_),
    .Q(\core.cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16006_ (.CLK(clk),
    .D(_00857_),
    .Q(\core.cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16007_ (.CLK(clk),
    .D(_00858_),
    .Q(\core.cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16008_ (.CLK(clk),
    .D(_00859_),
    .Q(\core.cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16009_ (.CLK(clk),
    .D(_00860_),
    .Q(\core.cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16010_ (.CLK(clk),
    .D(_00861_),
    .Q(\core.cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16011_ (.CLK(clk),
    .D(_00862_),
    .Q(\core.cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16012_ (.CLK(clk),
    .D(_00863_),
    .Q(\core.cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16013_ (.CLK(clk),
    .D(_00864_),
    .Q(\core.cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16014_ (.CLK(clk),
    .D(_00865_),
    .Q(\core.cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16015_ (.CLK(clk),
    .D(_00866_),
    .Q(\core.cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16016_ (.CLK(clk),
    .D(_00867_),
    .Q(\core.cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16017_ (.CLK(clk),
    .D(_00868_),
    .Q(\core.cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16018_ (.CLK(clk),
    .D(_00869_),
    .Q(\core.cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16019_ (.CLK(clk),
    .D(_00870_),
    .Q(\core.cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16020_ (.CLK(clk),
    .D(_00871_),
    .Q(\core.cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16021_ (.CLK(clk),
    .D(_00872_),
    .Q(\core.cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16022_ (.CLK(clk),
    .D(_00873_),
    .Q(\core.cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16023_ (.CLK(clk),
    .D(_00874_),
    .Q(\core.cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16024_ (.CLK(clk),
    .D(_00875_),
    .Q(\core.cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16025_ (.CLK(clk),
    .D(_00876_),
    .Q(\core.cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16026_ (.CLK(clk),
    .D(_00877_),
    .Q(\core.cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16027_ (.CLK(clk),
    .D(_00878_),
    .Q(\core.cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16028_ (.CLK(clk),
    .D(_00879_),
    .Q(\core.cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16029_ (.CLK(clk),
    .D(_00880_),
    .Q(\core.cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16030_ (.CLK(clk),
    .D(_00881_),
    .Q(\core.cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16031_ (.CLK(clk),
    .D(_00882_),
    .Q(\core.cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16032_ (.CLK(clk),
    .D(_00883_),
    .Q(\core.cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16033_ (.CLK(clk),
    .D(_00884_),
    .Q(\core.cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16034_ (.CLK(clk),
    .D(_00885_),
    .Q(\core.cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16035_ (.CLK(clk),
    .D(_00886_),
    .Q(\core.cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16036_ (.CLK(clk),
    .D(_00887_),
    .Q(\core.cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16037_ (.CLK(clk),
    .D(_00888_),
    .Q(\core.cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16038_ (.CLK(clk),
    .D(_00889_),
    .Q(\core.cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16039_ (.CLK(clk),
    .D(_00890_),
    .Q(\core.cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16040_ (.CLK(clk),
    .D(_00891_),
    .Q(\core.cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16041_ (.CLK(clk),
    .D(_00892_),
    .Q(\core.cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16042_ (.CLK(clk),
    .D(_00893_),
    .Q(\core.cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16043_ (.CLK(clk),
    .D(_00894_),
    .Q(\core.cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16044_ (.CLK(clk),
    .D(_00895_),
    .Q(\core.cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16045_ (.CLK(clk),
    .D(_00896_),
    .Q(\core.cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16046_ (.CLK(clk),
    .D(_00897_),
    .Q(\core.cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16047_ (.CLK(clk),
    .D(_00898_),
    .Q(\core.cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16048_ (.CLK(clk),
    .D(_00899_),
    .Q(\core.cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16049_ (.CLK(clk),
    .D(_00900_),
    .Q(\core.cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16050_ (.CLK(clk),
    .D(_00901_),
    .Q(\core.cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16051_ (.CLK(clk),
    .D(_00902_),
    .Q(\core.cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16052_ (.CLK(clk),
    .D(_00903_),
    .Q(\core.cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16053_ (.CLK(clk),
    .D(_00904_),
    .Q(\core.cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16054_ (.CLK(clk),
    .D(_00905_),
    .Q(\core.cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16055_ (.CLK(clk),
    .D(_00906_),
    .Q(\core.cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16056_ (.CLK(clk),
    .D(_00907_),
    .Q(\core.cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16057_ (.CLK(clk),
    .D(_00908_),
    .Q(\core.cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16058_ (.CLK(clk),
    .D(_00909_),
    .Q(\core.cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16059_ (.CLK(clk),
    .D(_00910_),
    .Q(\core.cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16060_ (.CLK(clk),
    .D(_00911_),
    .Q(\core.cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16061_ (.CLK(clk),
    .D(_00912_),
    .Q(\core.cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16062_ (.CLK(clk),
    .D(_00913_),
    .Q(\core.cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16063_ (.CLK(clk),
    .D(_00914_),
    .Q(\core.cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16064_ (.CLK(clk),
    .D(_00915_),
    .Q(\core.cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16065_ (.CLK(clk),
    .D(_00916_),
    .Q(\core.cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16066_ (.CLK(clk),
    .D(_00917_),
    .Q(\core.cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16067_ (.CLK(clk),
    .D(_00918_),
    .Q(\core.cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16068_ (.CLK(clk),
    .D(_00919_),
    .Q(\core.cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16069_ (.CLK(clk),
    .D(_00920_),
    .Q(\core.cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16070_ (.CLK(clk),
    .D(_00921_),
    .Q(\core.cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16071_ (.CLK(clk),
    .D(_00922_),
    .Q(\core.cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16072_ (.CLK(clk),
    .D(_00923_),
    .Q(\core.cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16073_ (.CLK(clk),
    .D(_00924_),
    .Q(\core.cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16074_ (.CLK(clk),
    .D(_00925_),
    .Q(\core.cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16075_ (.CLK(clk),
    .D(_00926_),
    .Q(\core.cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16076_ (.CLK(clk),
    .D(_00927_),
    .Q(\core.cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16077_ (.CLK(clk),
    .D(_00928_),
    .Q(\core.cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16078_ (.CLK(clk),
    .D(_00929_),
    .Q(\core.cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16079_ (.CLK(clk),
    .D(_00930_),
    .Q(\core.cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16080_ (.CLK(clk),
    .D(_00931_),
    .Q(\core.cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16081_ (.CLK(clk),
    .D(_00932_),
    .Q(\core.cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16082_ (.CLK(clk),
    .D(_00933_),
    .Q(\core.cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16083_ (.CLK(clk),
    .D(_00934_),
    .Q(\core.cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16084_ (.CLK(clk),
    .D(_00935_),
    .Q(\core.cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16085_ (.CLK(clk),
    .D(_00936_),
    .Q(\core.cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16086_ (.CLK(clk),
    .D(_00937_),
    .Q(\core.cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16087_ (.CLK(clk),
    .D(_00938_),
    .Q(\core.cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16088_ (.CLK(clk),
    .D(_00939_),
    .Q(\core.cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16089_ (.CLK(clk),
    .D(_00940_),
    .Q(\core.cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16090_ (.CLK(clk),
    .D(_00941_),
    .Q(\core.cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16091_ (.CLK(clk),
    .D(_00942_),
    .Q(\core.cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16092_ (.CLK(clk),
    .D(_00943_),
    .Q(\core.cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16093_ (.CLK(clk),
    .D(_00944_),
    .Q(\core.cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16094_ (.CLK(clk),
    .D(_00945_),
    .Q(\core.cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16095_ (.CLK(clk),
    .D(_00946_),
    .Q(\core.cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16096_ (.CLK(clk),
    .D(_00947_),
    .Q(\core.cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16097_ (.CLK(clk),
    .D(_00948_),
    .Q(\core.cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16098_ (.CLK(clk),
    .D(_00949_),
    .Q(\core.cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16099_ (.CLK(clk),
    .D(_00950_),
    .Q(\core.cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16100_ (.CLK(clk),
    .D(_00951_),
    .Q(\core.cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16101_ (.CLK(clk),
    .D(_00952_),
    .Q(\core.cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16102_ (.CLK(clk),
    .D(_00953_),
    .Q(\core.cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16103_ (.CLK(clk),
    .D(_00954_),
    .Q(\core.cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16104_ (.CLK(clk),
    .D(_00955_),
    .Q(\core.cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16105_ (.CLK(clk),
    .D(_00956_),
    .Q(\core.cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16106_ (.CLK(clk),
    .D(_00957_),
    .Q(\core.cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16107_ (.CLK(clk),
    .D(_00958_),
    .Q(\core.cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16108_ (.CLK(clk),
    .D(_00959_),
    .Q(\core.cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16109_ (.CLK(clk),
    .D(_00960_),
    .Q(\core.cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16110_ (.CLK(clk),
    .D(_00961_),
    .Q(\core.cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16111_ (.CLK(clk),
    .D(_00962_),
    .Q(\core.cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16112_ (.CLK(clk),
    .D(_00963_),
    .Q(\core.cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16113_ (.CLK(clk),
    .D(_00964_),
    .Q(\core.cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16114_ (.CLK(clk),
    .D(_00965_),
    .Q(\core.cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16115_ (.CLK(clk),
    .D(_00966_),
    .Q(\core.cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16116_ (.CLK(clk),
    .D(_00967_),
    .Q(\core.cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16117_ (.CLK(clk),
    .D(_00968_),
    .Q(\core.cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16118_ (.CLK(clk),
    .D(_00969_),
    .Q(\core.cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16119_ (.CLK(clk),
    .D(_00970_),
    .Q(\core.cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16120_ (.CLK(clk),
    .D(_00971_),
    .Q(\core.cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16121_ (.CLK(clk),
    .D(_00972_),
    .Q(\core.cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16122_ (.CLK(clk),
    .D(_00973_),
    .Q(\core.cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16123_ (.CLK(clk),
    .D(_00974_),
    .Q(\core.cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16124_ (.CLK(clk),
    .D(_00975_),
    .Q(\core.cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16125_ (.CLK(clk),
    .D(_00976_),
    .Q(\core.cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16126_ (.CLK(clk),
    .D(_00977_),
    .Q(\core.cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16127_ (.CLK(clk),
    .D(_00978_),
    .Q(\core.cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16128_ (.CLK(clk),
    .D(_00979_),
    .Q(\core.cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16129_ (.CLK(clk),
    .D(_00980_),
    .Q(\core.cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16130_ (.CLK(clk),
    .D(_00981_),
    .Q(\core.cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16131_ (.CLK(clk),
    .D(_00982_),
    .Q(\core.cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16132_ (.CLK(clk),
    .D(_00983_),
    .Q(\core.cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16133_ (.CLK(clk),
    .D(_00984_),
    .Q(\core.cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16134_ (.CLK(clk),
    .D(_00985_),
    .Q(\core.cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16135_ (.CLK(clk),
    .D(_00986_),
    .Q(\core.cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16136_ (.CLK(clk),
    .D(_00987_),
    .Q(\core.cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16137_ (.CLK(clk),
    .D(_00988_),
    .Q(\core.cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16138_ (.CLK(clk),
    .D(_00989_),
    .Q(\core.cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16139_ (.CLK(clk),
    .D(_00990_),
    .Q(\core.cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16140_ (.CLK(clk),
    .D(_00991_),
    .Q(\core.cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16141_ (.CLK(clk),
    .D(_00992_),
    .Q(\core.cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16142_ (.CLK(clk),
    .D(_00993_),
    .Q(\core.cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16143_ (.CLK(clk),
    .D(_00994_),
    .Q(\core.cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16144_ (.CLK(clk),
    .D(_00995_),
    .Q(\core.cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16145_ (.CLK(clk),
    .D(_00996_),
    .Q(\core.cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16146_ (.CLK(clk),
    .D(_00997_),
    .Q(\core.cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16147_ (.CLK(clk),
    .D(_00998_),
    .Q(\core.cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16148_ (.CLK(clk),
    .D(_00999_),
    .Q(\core.cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16149_ (.CLK(clk),
    .D(_01000_),
    .Q(\core.cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16150_ (.CLK(clk),
    .D(_01001_),
    .Q(\core.cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16151_ (.CLK(clk),
    .D(_01002_),
    .Q(\core.cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16152_ (.CLK(clk),
    .D(_01003_),
    .Q(\core.cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16153_ (.CLK(clk),
    .D(_01004_),
    .Q(\core.cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16154_ (.CLK(clk),
    .D(_01005_),
    .Q(\core.cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16155_ (.CLK(clk),
    .D(_01006_),
    .Q(\core.cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16156_ (.CLK(clk),
    .D(_01007_),
    .Q(\core.cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16157_ (.CLK(clk),
    .D(_01008_),
    .Q(\core.cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16158_ (.CLK(clk),
    .D(_01009_),
    .Q(\core.cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16159_ (.CLK(clk),
    .D(_01010_),
    .Q(\core.cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16160_ (.CLK(clk),
    .D(_01011_),
    .Q(\core.cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16161_ (.CLK(clk),
    .D(_01012_),
    .Q(\core.cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16162_ (.CLK(clk),
    .D(_01013_),
    .Q(\core.cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16163_ (.CLK(clk),
    .D(_01014_),
    .Q(\core.cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16164_ (.CLK(clk),
    .D(_01015_),
    .Q(\core.cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16165_ (.CLK(clk),
    .D(_01016_),
    .Q(\core.cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16166_ (.CLK(clk),
    .D(_01017_),
    .Q(\core.cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16167_ (.CLK(clk),
    .D(_01018_),
    .Q(\core.cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16168_ (.CLK(clk),
    .D(_01019_),
    .Q(\core.cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16169_ (.CLK(clk),
    .D(_01020_),
    .Q(\core.cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16170_ (.CLK(clk),
    .D(_01021_),
    .Q(\core.cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16171_ (.CLK(clk),
    .D(_01022_),
    .Q(\core.cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16172_ (.CLK(clk),
    .D(_01023_),
    .Q(\core.cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16173_ (.CLK(clk),
    .D(_01024_),
    .Q(\core.cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16174_ (.CLK(clk),
    .D(_01025_),
    .Q(\core.cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16175_ (.CLK(clk),
    .D(_01026_),
    .Q(\core.cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16176_ (.CLK(clk),
    .D(_01027_),
    .Q(\core.cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16177_ (.CLK(clk),
    .D(_01028_),
    .Q(\core.cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16178_ (.CLK(clk),
    .D(_01029_),
    .Q(\core.cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16179_ (.CLK(clk),
    .D(_01030_),
    .Q(\core.cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16180_ (.CLK(clk),
    .D(_01031_),
    .Q(\core.cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16181_ (.CLK(clk),
    .D(_01032_),
    .Q(\core.cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16182_ (.CLK(clk),
    .D(_01033_),
    .Q(\core.cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16183_ (.CLK(clk),
    .D(_01034_),
    .Q(\core.cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16184_ (.CLK(clk),
    .D(_01035_),
    .Q(\core.cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16185_ (.CLK(clk),
    .D(_01036_),
    .Q(\core.cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16186_ (.CLK(clk),
    .D(_01037_),
    .Q(\core.cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16187_ (.CLK(clk),
    .D(_01038_),
    .Q(\core.cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16188_ (.CLK(clk),
    .D(_01039_),
    .Q(\core.cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16189_ (.CLK(clk),
    .D(_01040_),
    .Q(\core.cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16190_ (.CLK(clk),
    .D(_01041_),
    .Q(\core.cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16191_ (.CLK(clk),
    .D(_01042_),
    .Q(\core.cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16192_ (.CLK(clk),
    .D(_01043_),
    .Q(\core.cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16193_ (.CLK(clk),
    .D(_01044_),
    .Q(\core.cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16194_ (.CLK(clk),
    .D(_01045_),
    .Q(\core.cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16195_ (.CLK(clk),
    .D(_01046_),
    .Q(\core.cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16196_ (.CLK(clk),
    .D(_01047_),
    .Q(\core.cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16197_ (.CLK(clk),
    .D(_01048_),
    .Q(\core.cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16198_ (.CLK(clk),
    .D(_01049_),
    .Q(\core.cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16199_ (.CLK(clk),
    .D(_01050_),
    .Q(\core.cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16200_ (.CLK(clk),
    .D(_01051_),
    .Q(\core.cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16201_ (.CLK(clk),
    .D(_01052_),
    .Q(\core.cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16202_ (.CLK(clk),
    .D(_01053_),
    .Q(\core.cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16203_ (.CLK(clk),
    .D(_01054_),
    .Q(\core.cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16204_ (.CLK(clk),
    .D(_01055_),
    .Q(\core.cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16205_ (.CLK(clk),
    .D(_01056_),
    .Q(\core.cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16206_ (.CLK(clk),
    .D(_01057_),
    .Q(\core.cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16207_ (.CLK(clk),
    .D(_01058_),
    .Q(\core.cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16208_ (.CLK(clk),
    .D(_01059_),
    .Q(\core.cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16209_ (.CLK(clk),
    .D(_01060_),
    .Q(\core.cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16210_ (.CLK(clk),
    .D(_01061_),
    .Q(\core.cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16211_ (.CLK(clk),
    .D(_01062_),
    .Q(\core.cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16212_ (.CLK(clk),
    .D(_01063_),
    .Q(\core.cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16213_ (.CLK(clk),
    .D(_01064_),
    .Q(\core.cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16214_ (.CLK(clk),
    .D(_01065_),
    .Q(\core.cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16215_ (.CLK(clk),
    .D(_01066_),
    .Q(\core.cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16216_ (.CLK(clk),
    .D(_01067_),
    .Q(\core.cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16217_ (.CLK(clk),
    .D(_01068_),
    .Q(\core.cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16218_ (.CLK(clk),
    .D(_01069_),
    .Q(\core.cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16219_ (.CLK(clk),
    .D(_01070_),
    .Q(\core.cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16220_ (.CLK(clk),
    .D(_01071_),
    .Q(\core.cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16221_ (.CLK(clk),
    .D(_01072_),
    .Q(\core.cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16222_ (.CLK(clk),
    .D(_01073_),
    .Q(\core.cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16223_ (.CLK(clk),
    .D(_01074_),
    .Q(\core.cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16224_ (.CLK(clk),
    .D(_01075_),
    .Q(\core.cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16225_ (.CLK(clk),
    .D(_01076_),
    .Q(\core.cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16226_ (.CLK(clk),
    .D(_01077_),
    .Q(\core.cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16227_ (.CLK(clk),
    .D(_01078_),
    .Q(\core.cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16228_ (.CLK(clk),
    .D(_01079_),
    .Q(\core.cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16229_ (.CLK(clk),
    .D(_01080_),
    .Q(\core.cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16230_ (.CLK(clk),
    .D(_01081_),
    .Q(\core.cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16231_ (.CLK(clk),
    .D(_01082_),
    .Q(\core.cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16232_ (.CLK(clk),
    .D(_01083_),
    .Q(\core.cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16233_ (.CLK(clk),
    .D(_01084_),
    .Q(\core.cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16234_ (.CLK(clk),
    .D(_01085_),
    .Q(\core.cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16235_ (.CLK(clk),
    .D(_01086_),
    .Q(\core.cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16236_ (.CLK(clk),
    .D(_01087_),
    .Q(\core.cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16237_ (.CLK(clk),
    .D(_01088_),
    .Q(\core.cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16238_ (.CLK(clk),
    .D(_01089_),
    .Q(\core.cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16239_ (.CLK(clk),
    .D(_01090_),
    .Q(\core.cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16240_ (.CLK(clk),
    .D(_01091_),
    .Q(\core.cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16241_ (.CLK(clk),
    .D(_01092_),
    .Q(\core.cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16242_ (.CLK(clk),
    .D(_01093_),
    .Q(\core.cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16243_ (.CLK(clk),
    .D(_01094_),
    .Q(\core.cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16244_ (.CLK(clk),
    .D(_01095_),
    .Q(\core.cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16245_ (.CLK(clk),
    .D(_01096_),
    .Q(\core.cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16246_ (.CLK(clk),
    .D(_01097_),
    .Q(\core.cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16247_ (.CLK(clk),
    .D(_01098_),
    .Q(\core.cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16248_ (.CLK(clk),
    .D(_01099_),
    .Q(\core.cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16249_ (.CLK(clk),
    .D(_01100_),
    .Q(\core.cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16250_ (.CLK(clk),
    .D(_01101_),
    .Q(\core.cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16251_ (.CLK(clk),
    .D(_01102_),
    .Q(\core.cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16252_ (.CLK(clk),
    .D(_01103_),
    .Q(\core.cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16253_ (.CLK(clk),
    .D(_01104_),
    .Q(\core.cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16254_ (.CLK(clk),
    .D(_01105_),
    .Q(\core.cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16255_ (.CLK(clk),
    .D(_01106_),
    .Q(\core.cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16256_ (.CLK(clk),
    .D(_01107_),
    .Q(\core.cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16257_ (.CLK(clk),
    .D(_01108_),
    .Q(\core.cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16258_ (.CLK(clk),
    .D(_01109_),
    .Q(\core.cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16259_ (.CLK(clk),
    .D(_01110_),
    .Q(\core.cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16260_ (.CLK(clk),
    .D(_01111_),
    .Q(\core.cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16261_ (.CLK(clk),
    .D(_01112_),
    .Q(\core.cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16262_ (.CLK(clk),
    .D(_01113_),
    .Q(\core.cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16263_ (.CLK(clk),
    .D(_01114_),
    .Q(\core.cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16264_ (.CLK(clk),
    .D(_01115_),
    .Q(\core.cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16265_ (.CLK(clk),
    .D(_01116_),
    .Q(\core.cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16266_ (.CLK(clk),
    .D(_01117_),
    .Q(\core.cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16267_ (.CLK(clk),
    .D(_01118_),
    .Q(\core.cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16268_ (.CLK(clk),
    .D(_01119_),
    .Q(\core.cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16269_ (.CLK(clk),
    .D(_01120_),
    .Q(\core.cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16270_ (.CLK(clk),
    .D(_01121_),
    .Q(\core.cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16271_ (.CLK(clk),
    .D(_01122_),
    .Q(\core.cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16272_ (.CLK(clk),
    .D(_01123_),
    .Q(\core.cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16273_ (.CLK(clk),
    .D(_01124_),
    .Q(\core.cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16274_ (.CLK(clk),
    .D(_01125_),
    .Q(\core.cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16275_ (.CLK(clk),
    .D(_01126_),
    .Q(\core.cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16276_ (.CLK(clk),
    .D(_01127_),
    .Q(\core.cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16277_ (.CLK(clk),
    .D(_01128_),
    .Q(\core.cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16278_ (.CLK(clk),
    .D(_01129_),
    .Q(\core.cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16279_ (.CLK(clk),
    .D(_01130_),
    .Q(\core.cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16280_ (.CLK(clk),
    .D(_01131_),
    .Q(\core.cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16281_ (.CLK(clk),
    .D(_01132_),
    .Q(\core.cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16282_ (.CLK(clk),
    .D(_01133_),
    .Q(\core.cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16283_ (.CLK(clk),
    .D(_01134_),
    .Q(\core.cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16284_ (.CLK(clk),
    .D(_01135_),
    .Q(\core.cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16285_ (.CLK(clk),
    .D(_01136_),
    .Q(\core.cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16286_ (.CLK(clk),
    .D(_01137_),
    .Q(\core.cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16287_ (.CLK(clk),
    .D(_01138_),
    .Q(\core.cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16288_ (.CLK(clk),
    .D(_01139_),
    .Q(\core.cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16289_ (.CLK(clk),
    .D(_01140_),
    .Q(\core.cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16290_ (.CLK(clk),
    .D(_01141_),
    .Q(\core.cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16291_ (.CLK(clk),
    .D(_01142_),
    .Q(\core.cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16292_ (.CLK(clk),
    .D(_01143_),
    .Q(\core.cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16293_ (.CLK(clk),
    .D(_01144_),
    .Q(\core.cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16294_ (.CLK(clk),
    .D(_01145_),
    .Q(\core.cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16295_ (.CLK(clk),
    .D(_01146_),
    .Q(\core.cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16296_ (.CLK(clk),
    .D(_01147_),
    .Q(\core.cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16297_ (.CLK(clk),
    .D(_01148_),
    .Q(\core.cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16298_ (.CLK(clk),
    .D(_01149_),
    .Q(\core.cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16299_ (.CLK(clk),
    .D(_01150_),
    .Q(\core.cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16300_ (.CLK(clk),
    .D(_01151_),
    .Q(\core.cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16301_ (.CLK(clk),
    .D(_01152_),
    .Q(\core.cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16302_ (.CLK(clk),
    .D(_01153_),
    .Q(\core.cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16303_ (.CLK(clk),
    .D(_01154_),
    .Q(\core.cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16304_ (.CLK(clk),
    .D(_01155_),
    .Q(\core.cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16305_ (.CLK(clk),
    .D(_01156_),
    .Q(\core.cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16306_ (.CLK(clk),
    .D(_01157_),
    .Q(\core.cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16307_ (.CLK(clk),
    .D(_01158_),
    .Q(\core.cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16308_ (.CLK(clk),
    .D(_01159_),
    .Q(\core.cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16309_ (.CLK(clk),
    .D(_01160_),
    .Q(\core.cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16310_ (.CLK(clk),
    .D(_01161_),
    .Q(\core.cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16311_ (.CLK(clk),
    .D(_01162_),
    .Q(\core.cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16312_ (.CLK(clk),
    .D(_01163_),
    .Q(\core.cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16313_ (.CLK(clk),
    .D(_01164_),
    .Q(\core.cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16314_ (.CLK(clk),
    .D(_01165_),
    .Q(\core.cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16315_ (.CLK(clk),
    .D(_01166_),
    .Q(\core.cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16316_ (.CLK(clk),
    .D(_01167_),
    .Q(\core.cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16317_ (.CLK(clk),
    .D(_01168_),
    .Q(\core.cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16318_ (.CLK(clk),
    .D(_01169_),
    .Q(\core.cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16319_ (.CLK(clk),
    .D(_01170_),
    .Q(\core.cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16320_ (.CLK(clk),
    .D(_01171_),
    .Q(\core.cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16321_ (.CLK(clk),
    .D(_01172_),
    .Q(\core.cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16322_ (.CLK(clk),
    .D(_01173_),
    .Q(\core.cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16323_ (.CLK(clk),
    .D(_01174_),
    .Q(\core.cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16324_ (.CLK(clk),
    .D(_01175_),
    .Q(\core.cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16325_ (.CLK(clk),
    .D(_01176_),
    .Q(\core.cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16326_ (.CLK(clk),
    .D(_01177_),
    .Q(\core.cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16327_ (.CLK(clk),
    .D(_01178_),
    .Q(\core.cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16328_ (.CLK(clk),
    .D(_01179_),
    .Q(\core.cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16329_ (.CLK(clk),
    .D(_01180_),
    .Q(\core.cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16330_ (.CLK(clk),
    .D(_01181_),
    .Q(\core.cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16331_ (.CLK(clk),
    .D(_01182_),
    .Q(\core.cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16332_ (.CLK(clk),
    .D(_01183_),
    .Q(\core.cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16333_ (.CLK(clk),
    .D(_01184_),
    .Q(\core.cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16334_ (.CLK(clk),
    .D(_01185_),
    .Q(\core.cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16335_ (.CLK(clk),
    .D(_01186_),
    .Q(\core.cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16336_ (.CLK(clk),
    .D(_01187_),
    .Q(\core.cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16337_ (.CLK(clk),
    .D(_01188_),
    .Q(\core.cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16338_ (.CLK(clk),
    .D(_01189_),
    .Q(\core.cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16339_ (.CLK(clk),
    .D(_01190_),
    .Q(\core.cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16340_ (.CLK(clk),
    .D(_01191_),
    .Q(\core.cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16341_ (.CLK(clk),
    .D(_01192_),
    .Q(\core.cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16342_ (.CLK(clk),
    .D(_01193_),
    .Q(\core.cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16343_ (.CLK(clk),
    .D(_01194_),
    .Q(\core.cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16344_ (.CLK(clk),
    .D(_01195_),
    .Q(\core.cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16345_ (.CLK(clk),
    .D(_01196_),
    .Q(\core.cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16346_ (.CLK(clk),
    .D(_01197_),
    .Q(\core.cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16347_ (.CLK(clk),
    .D(_01198_),
    .Q(\core.cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16348_ (.CLK(clk),
    .D(_01199_),
    .Q(\core.cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16349_ (.CLK(clk),
    .D(_01200_),
    .Q(\core.cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16350_ (.CLK(clk),
    .D(_01201_),
    .Q(\core.cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16351_ (.CLK(clk),
    .D(_01202_),
    .Q(\core.cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16352_ (.CLK(clk),
    .D(_01203_),
    .Q(\core.cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16353_ (.CLK(clk),
    .D(_01204_),
    .Q(\core.cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16354_ (.CLK(clk),
    .D(_01205_),
    .Q(\core.cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16355_ (.CLK(clk),
    .D(_01206_),
    .Q(\core.cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16356_ (.CLK(clk),
    .D(_01207_),
    .Q(\core.cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16357_ (.CLK(clk),
    .D(_01208_),
    .Q(\core.cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16358_ (.CLK(clk),
    .D(_01209_),
    .Q(\core.cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16359_ (.CLK(clk),
    .D(_01210_),
    .Q(\core.cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16360_ (.CLK(clk),
    .D(_01211_),
    .Q(\core.cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16361_ (.CLK(clk),
    .D(_01212_),
    .Q(\core.cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16362_ (.CLK(clk),
    .D(_01213_),
    .Q(\core.cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16363_ (.CLK(clk),
    .D(_01214_),
    .Q(\core.cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16364_ (.CLK(clk),
    .D(_01215_),
    .Q(\core.cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16365_ (.CLK(clk),
    .D(_01216_),
    .Q(\core.cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16366_ (.CLK(clk),
    .D(_01217_),
    .Q(\core.cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16367_ (.CLK(clk),
    .D(_01218_),
    .Q(\core.cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16368_ (.CLK(clk),
    .D(_01219_),
    .Q(\core.cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16369_ (.CLK(clk),
    .D(_01220_),
    .Q(\core.cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16370_ (.CLK(clk),
    .D(_01221_),
    .Q(\core.cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16371_ (.CLK(clk),
    .D(_01222_),
    .Q(\core.cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16372_ (.CLK(clk),
    .D(_01223_),
    .Q(\core.cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16373_ (.CLK(clk),
    .D(_01224_),
    .Q(\core.cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16374_ (.CLK(clk),
    .D(_01225_),
    .Q(\core.cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16375_ (.CLK(clk),
    .D(_01226_),
    .Q(\core.cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16376_ (.CLK(clk),
    .D(_01227_),
    .Q(\core.cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16377_ (.CLK(clk),
    .D(_01228_),
    .Q(\core.cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16378_ (.CLK(clk),
    .D(_01229_),
    .Q(\core.cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16379_ (.CLK(clk),
    .D(_01230_),
    .Q(\core.cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16380_ (.CLK(clk),
    .D(_01231_),
    .Q(\core.cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16381_ (.CLK(clk),
    .D(_01232_),
    .Q(\core.cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16382_ (.CLK(clk),
    .D(_01233_),
    .Q(\core.cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16383_ (.CLK(clk),
    .D(_01234_),
    .Q(\core.cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16384_ (.CLK(clk),
    .D(_01235_),
    .Q(\core.cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16385_ (.CLK(clk),
    .D(_01236_),
    .Q(\core.cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16386_ (.CLK(clk),
    .D(_01237_),
    .Q(\core.cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16387_ (.CLK(clk),
    .D(_01238_),
    .Q(\core.cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16388_ (.CLK(clk),
    .D(_01239_),
    .Q(\core.cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16389_ (.CLK(clk),
    .D(_01240_),
    .Q(\core.cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16390_ (.CLK(clk),
    .D(_01241_),
    .Q(\core.cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16391_ (.CLK(clk),
    .D(_01242_),
    .Q(\core.cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16392_ (.CLK(clk),
    .D(_01243_),
    .Q(\core.cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16393_ (.CLK(clk),
    .D(_01244_),
    .Q(\core.cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16394_ (.CLK(clk),
    .D(_01245_),
    .Q(\core.cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16395_ (.CLK(clk),
    .D(_01246_),
    .Q(\core.cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16396_ (.CLK(clk),
    .D(_00017_),
    .Q(\core.mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_2 _16397_ (.CLK(clk),
    .D(_00018_),
    .Q(\core.mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16398_ (.CLK(clk),
    .D(_00019_),
    .Q(\core.mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_2 _16399_ (.CLK(clk),
    .D(_01247_),
    .Q(\core.cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16400_ (.CLK(clk),
    .D(_01248_),
    .Q(\core.cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16401_ (.CLK(clk),
    .D(_01249_),
    .Q(\core.cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16402_ (.CLK(clk),
    .D(_01250_),
    .Q(\core.cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16403_ (.CLK(clk),
    .D(_01251_),
    .Q(\core.cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16404_ (.CLK(clk),
    .D(_01252_),
    .Q(\core.cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16405_ (.CLK(clk),
    .D(_01253_),
    .Q(\core.cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16406_ (.CLK(clk),
    .D(_01254_),
    .Q(\core.cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16407_ (.CLK(clk),
    .D(_01255_),
    .Q(\core.cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16408_ (.CLK(clk),
    .D(_01256_),
    .Q(\core.cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16409_ (.CLK(clk),
    .D(_01257_),
    .Q(\core.cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16410_ (.CLK(clk),
    .D(_01258_),
    .Q(\core.cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16411_ (.CLK(clk),
    .D(_01259_),
    .Q(\core.cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16412_ (.CLK(clk),
    .D(_01260_),
    .Q(\core.cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16413_ (.CLK(clk),
    .D(_01261_),
    .Q(\core.cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16414_ (.CLK(clk),
    .D(_01262_),
    .Q(\core.cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16415_ (.CLK(clk),
    .D(_01263_),
    .Q(\core.cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16416_ (.CLK(clk),
    .D(_01264_),
    .Q(\core.cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16417_ (.CLK(clk),
    .D(_01265_),
    .Q(\core.cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16418_ (.CLK(clk),
    .D(_01266_),
    .Q(\core.cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16419_ (.CLK(clk),
    .D(_01267_),
    .Q(\core.cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16420_ (.CLK(clk),
    .D(_01268_),
    .Q(\core.cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16421_ (.CLK(clk),
    .D(_01269_),
    .Q(\core.cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16422_ (.CLK(clk),
    .D(_01270_),
    .Q(\core.cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16423_ (.CLK(clk),
    .D(_01271_),
    .Q(\core.cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16424_ (.CLK(clk),
    .D(_01272_),
    .Q(\core.cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16425_ (.CLK(clk),
    .D(_01273_),
    .Q(\core.cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16426_ (.CLK(clk),
    .D(_01274_),
    .Q(\core.cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16427_ (.CLK(clk),
    .D(_01275_),
    .Q(\core.cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16428_ (.CLK(clk),
    .D(_01276_),
    .Q(\core.cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16429_ (.CLK(clk),
    .D(_01277_),
    .Q(\core.cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16430_ (.CLK(clk),
    .D(_01278_),
    .Q(\core.cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16431_ (.CLK(clk),
    .D(_00010_),
    .Q(\core.cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _16432_ (.CLK(clk),
    .D(_00011_),
    .Q(\core.cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16433_ (.CLK(clk),
    .D(_00012_),
    .Q(\core.cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _16434_ (.CLK(clk),
    .D(_00013_),
    .Q(\core.cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _16435_ (.CLK(clk),
    .D(_00014_),
    .Q(\core.cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _16436_ (.CLK(clk),
    .D(_00015_),
    .Q(\core.cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _16437_ (.CLK(clk),
    .D(_00016_),
    .Q(\core.cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_2 _16438_ (.CLK(clk),
    .D(_01279_),
    .Q(\core.cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16439_ (.CLK(clk),
    .D(_01280_),
    .Q(\core.cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16440_ (.CLK(clk),
    .D(_01281_),
    .Q(\core.cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16441_ (.CLK(clk),
    .D(_01282_),
    .Q(\core.cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16442_ (.CLK(clk),
    .D(_01283_),
    .Q(\core.cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16443_ (.CLK(clk),
    .D(_01284_),
    .Q(\core.cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16444_ (.CLK(clk),
    .D(_01285_),
    .Q(\core.cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16445_ (.CLK(clk),
    .D(_01286_),
    .Q(\core.cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16446_ (.CLK(clk),
    .D(_01287_),
    .Q(\core.cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16447_ (.CLK(clk),
    .D(_01288_),
    .Q(\core.cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16448_ (.CLK(clk),
    .D(_01289_),
    .Q(\core.cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16449_ (.CLK(clk),
    .D(_01290_),
    .Q(\core.cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16450_ (.CLK(clk),
    .D(_01291_),
    .Q(\core.cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16451_ (.CLK(clk),
    .D(_01292_),
    .Q(\core.cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16452_ (.CLK(clk),
    .D(_01293_),
    .Q(\core.cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16453_ (.CLK(clk),
    .D(_01294_),
    .Q(\core.cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16454_ (.CLK(clk),
    .D(_01295_),
    .Q(\core.cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16455_ (.CLK(clk),
    .D(_01296_),
    .Q(\core.cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16456_ (.CLK(clk),
    .D(_01297_),
    .Q(\core.cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16457_ (.CLK(clk),
    .D(_01298_),
    .Q(\core.cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16458_ (.CLK(clk),
    .D(_01299_),
    .Q(\core.cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16459_ (.CLK(clk),
    .D(_01300_),
    .Q(\core.cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16460_ (.CLK(clk),
    .D(_01301_),
    .Q(\core.cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16461_ (.CLK(clk),
    .D(_01302_),
    .Q(\core.cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16462_ (.CLK(clk),
    .D(_01303_),
    .Q(\core.cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16463_ (.CLK(clk),
    .D(_01304_),
    .Q(\core.cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16464_ (.CLK(clk),
    .D(_01305_),
    .Q(\core.cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16465_ (.CLK(clk),
    .D(_01306_),
    .Q(\core.cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16466_ (.CLK(clk),
    .D(_01307_),
    .Q(\core.cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16467_ (.CLK(clk),
    .D(_01308_),
    .Q(\core.cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16468_ (.CLK(clk),
    .D(_01309_),
    .Q(\core.cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16469_ (.CLK(clk),
    .D(_01310_),
    .Q(\core.cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16470_ (.CLK(clk),
    .D(_01311_),
    .Q(\core.cpuregs[31][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16471_ (.CLK(clk),
    .D(_01312_),
    .Q(\core.cpuregs[31][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16472_ (.CLK(clk),
    .D(_01313_),
    .Q(\core.cpuregs[31][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16473_ (.CLK(clk),
    .D(_01314_),
    .Q(\core.cpuregs[31][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16474_ (.CLK(clk),
    .D(_01315_),
    .Q(\core.cpuregs[31][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16475_ (.CLK(clk),
    .D(_01316_),
    .Q(\core.cpuregs[31][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16476_ (.CLK(clk),
    .D(_01317_),
    .Q(\core.cpuregs[31][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16477_ (.CLK(clk),
    .D(_01318_),
    .Q(\core.cpuregs[31][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16478_ (.CLK(clk),
    .D(_01319_),
    .Q(\core.cpuregs[31][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16479_ (.CLK(clk),
    .D(_01320_),
    .Q(\core.cpuregs[31][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16480_ (.CLK(clk),
    .D(_01321_),
    .Q(\core.cpuregs[31][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16481_ (.CLK(clk),
    .D(_01322_),
    .Q(\core.cpuregs[31][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16482_ (.CLK(clk),
    .D(_01323_),
    .Q(\core.cpuregs[31][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16483_ (.CLK(clk),
    .D(_01324_),
    .Q(\core.cpuregs[31][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16484_ (.CLK(clk),
    .D(_01325_),
    .Q(\core.cpuregs[31][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16485_ (.CLK(clk),
    .D(_01326_),
    .Q(\core.cpuregs[31][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16486_ (.CLK(clk),
    .D(_01327_),
    .Q(\core.cpuregs[31][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16487_ (.CLK(clk),
    .D(_01328_),
    .Q(\core.cpuregs[31][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16488_ (.CLK(clk),
    .D(_01329_),
    .Q(\core.cpuregs[31][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16489_ (.CLK(clk),
    .D(_01330_),
    .Q(\core.cpuregs[31][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16490_ (.CLK(clk),
    .D(_01331_),
    .Q(\core.cpuregs[31][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16491_ (.CLK(clk),
    .D(_01332_),
    .Q(\core.cpuregs[31][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16492_ (.CLK(clk),
    .D(_01333_),
    .Q(\core.cpuregs[31][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16493_ (.CLK(clk),
    .D(_01334_),
    .Q(\core.cpuregs[31][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16494_ (.CLK(clk),
    .D(_01335_),
    .Q(\core.cpuregs[31][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16495_ (.CLK(clk),
    .D(_01336_),
    .Q(\core.cpuregs[31][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16496_ (.CLK(clk),
    .D(_01337_),
    .Q(\core.cpuregs[31][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16497_ (.CLK(clk),
    .D(_01338_),
    .Q(\core.cpuregs[31][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16498_ (.CLK(clk),
    .D(_01339_),
    .Q(\core.cpuregs[31][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16499_ (.CLK(clk),
    .D(_01340_),
    .Q(\core.cpuregs[31][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16500_ (.CLK(clk),
    .D(_01341_),
    .Q(\core.cpuregs[31][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16501_ (.CLK(clk),
    .D(_01342_),
    .Q(\core.cpuregs[31][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16502_ (.CLK(clk),
    .D(_01343_),
    .Q(\core.mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _16503_ (.CLK(clk),
    .D(_01344_),
    .Q(\core.mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16504_ (.CLK(clk),
    .D(_01345_),
    .Q(\core.mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _16505_ (.CLK(clk),
    .D(_01346_),
    .Q(\core.mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _16506_ (.CLK(clk),
    .D(_01347_),
    .Q(\core.mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _16507_ (.CLK(clk),
    .D(_01348_),
    .Q(\core.mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _16508_ (.CLK(clk),
    .D(_01349_),
    .Q(\core.mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _16509_ (.CLK(clk),
    .D(_01350_),
    .Q(\core.mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _16510_ (.CLK(clk),
    .D(_01351_),
    .Q(\core.mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _16511_ (.CLK(clk),
    .D(_01352_),
    .Q(\core.mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _16512_ (.CLK(clk),
    .D(_01353_),
    .Q(\core.mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _16513_ (.CLK(clk),
    .D(_01354_),
    .Q(\core.mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _16514_ (.CLK(clk),
    .D(_01355_),
    .Q(\core.mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _16515_ (.CLK(clk),
    .D(_01356_),
    .Q(\core.mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _16516_ (.CLK(clk),
    .D(_01357_),
    .Q(\core.mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _16517_ (.CLK(clk),
    .D(_01358_),
    .Q(\core.mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _16518_ (.CLK(clk),
    .D(_01359_),
    .Q(\core.mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _16519_ (.CLK(clk),
    .D(_01360_),
    .Q(\core.mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _16520_ (.CLK(clk),
    .D(_01361_),
    .Q(\core.mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _16521_ (.CLK(clk),
    .D(_01362_),
    .Q(\core.mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _16522_ (.CLK(clk),
    .D(_01363_),
    .Q(\core.mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _16523_ (.CLK(clk),
    .D(_01364_),
    .Q(\core.mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _16524_ (.CLK(clk),
    .D(_01365_),
    .Q(\core.mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _16525_ (.CLK(clk),
    .D(_01366_),
    .Q(\core.mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _16526_ (.CLK(clk),
    .D(_01367_),
    .Q(\core.mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _16527_ (.CLK(clk),
    .D(_01368_),
    .Q(\core.mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _16528_ (.CLK(clk),
    .D(_01369_),
    .Q(\core.mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _16529_ (.CLK(clk),
    .D(_01370_),
    .Q(\core.mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _16530_ (.CLK(clk),
    .D(_01371_),
    .Q(\core.mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _16531_ (.CLK(clk),
    .D(_01372_),
    .Q(\core.mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _16532_ (.CLK(clk),
    .D(_01373_),
    .Q(\core.mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _16533_ (.CLK(clk),
    .D(_01374_),
    .Q(\core.mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _16534_ (.CLK(clk),
    .D(_00025_),
    .Q(_00005_));
 sky130_fd_sc_hd__dfxtp_2 _16535_ (.CLK(clk),
    .D(_00026_),
    .Q(_00006_));
 sky130_fd_sc_hd__dfxtp_2 _16536_ (.CLK(clk),
    .D(_00027_),
    .Q(_00007_));
 sky130_fd_sc_hd__dfxtp_2 _16537_ (.CLK(clk),
    .D(_00028_),
    .Q(_00008_));
 sky130_fd_sc_hd__dfxtp_2 _16538_ (.CLK(clk),
    .D(_00029_),
    .Q(_00009_));
 sky130_fd_sc_hd__dfxtp_2 _16539_ (.CLK(clk),
    .D(_01375_),
    .Q(\core.cpuregs[29][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16540_ (.CLK(clk),
    .D(_01376_),
    .Q(\core.cpuregs[29][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16541_ (.CLK(clk),
    .D(_01377_),
    .Q(\core.cpuregs[29][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16542_ (.CLK(clk),
    .D(_01378_),
    .Q(\core.cpuregs[29][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16543_ (.CLK(clk),
    .D(_01379_),
    .Q(\core.cpuregs[29][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16544_ (.CLK(clk),
    .D(_01380_),
    .Q(\core.cpuregs[29][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16545_ (.CLK(clk),
    .D(_01381_),
    .Q(\core.cpuregs[29][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16546_ (.CLK(clk),
    .D(_01382_),
    .Q(\core.cpuregs[29][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16547_ (.CLK(clk),
    .D(_01383_),
    .Q(\core.cpuregs[29][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16548_ (.CLK(clk),
    .D(_01384_),
    .Q(\core.cpuregs[29][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16549_ (.CLK(clk),
    .D(_01385_),
    .Q(\core.cpuregs[29][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16550_ (.CLK(clk),
    .D(_01386_),
    .Q(\core.cpuregs[29][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16551_ (.CLK(clk),
    .D(_01387_),
    .Q(\core.cpuregs[29][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16552_ (.CLK(clk),
    .D(_01388_),
    .Q(\core.cpuregs[29][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16553_ (.CLK(clk),
    .D(_01389_),
    .Q(\core.cpuregs[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16554_ (.CLK(clk),
    .D(_01390_),
    .Q(\core.cpuregs[29][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16555_ (.CLK(clk),
    .D(_01391_),
    .Q(\core.cpuregs[29][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16556_ (.CLK(clk),
    .D(_01392_),
    .Q(\core.cpuregs[29][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16557_ (.CLK(clk),
    .D(_01393_),
    .Q(\core.cpuregs[29][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16558_ (.CLK(clk),
    .D(_01394_),
    .Q(\core.cpuregs[29][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16559_ (.CLK(clk),
    .D(_01395_),
    .Q(\core.cpuregs[29][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16560_ (.CLK(clk),
    .D(_01396_),
    .Q(\core.cpuregs[29][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16561_ (.CLK(clk),
    .D(_01397_),
    .Q(\core.cpuregs[29][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16562_ (.CLK(clk),
    .D(_01398_),
    .Q(\core.cpuregs[29][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16563_ (.CLK(clk),
    .D(_01399_),
    .Q(\core.cpuregs[29][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16564_ (.CLK(clk),
    .D(_01400_),
    .Q(\core.cpuregs[29][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16565_ (.CLK(clk),
    .D(_01401_),
    .Q(\core.cpuregs[29][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16566_ (.CLK(clk),
    .D(_01402_),
    .Q(\core.cpuregs[29][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16567_ (.CLK(clk),
    .D(_01403_),
    .Q(\core.cpuregs[29][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16568_ (.CLK(clk),
    .D(_01404_),
    .Q(\core.cpuregs[29][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16569_ (.CLK(clk),
    .D(_01405_),
    .Q(\core.cpuregs[29][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16570_ (.CLK(clk),
    .D(_01406_),
    .Q(\core.cpuregs[29][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16571_ (.CLK(clk),
    .D(_01407_),
    .Q(\core.cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16572_ (.CLK(clk),
    .D(_01408_),
    .Q(\core.cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16573_ (.CLK(clk),
    .D(_01409_),
    .Q(\core.cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16574_ (.CLK(clk),
    .D(_01410_),
    .Q(\core.cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16575_ (.CLK(clk),
    .D(_01411_),
    .Q(\core.cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16576_ (.CLK(clk),
    .D(_01412_),
    .Q(\core.cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16577_ (.CLK(clk),
    .D(_01413_),
    .Q(\core.cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16578_ (.CLK(clk),
    .D(_01414_),
    .Q(\core.cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16579_ (.CLK(clk),
    .D(_01415_),
    .Q(\core.cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16580_ (.CLK(clk),
    .D(_01416_),
    .Q(\core.cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16581_ (.CLK(clk),
    .D(_01417_),
    .Q(\core.cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16582_ (.CLK(clk),
    .D(_01418_),
    .Q(\core.cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16583_ (.CLK(clk),
    .D(_01419_),
    .Q(\core.cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16584_ (.CLK(clk),
    .D(_01420_),
    .Q(\core.cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16585_ (.CLK(clk),
    .D(_01421_),
    .Q(\core.cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16586_ (.CLK(clk),
    .D(_01422_),
    .Q(\core.cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16587_ (.CLK(clk),
    .D(_01423_),
    .Q(\core.cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16588_ (.CLK(clk),
    .D(_01424_),
    .Q(\core.cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16589_ (.CLK(clk),
    .D(_01425_),
    .Q(\core.cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16590_ (.CLK(clk),
    .D(_01426_),
    .Q(\core.cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16591_ (.CLK(clk),
    .D(_01427_),
    .Q(\core.cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16592_ (.CLK(clk),
    .D(_01428_),
    .Q(\core.cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16593_ (.CLK(clk),
    .D(_01429_),
    .Q(\core.cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16594_ (.CLK(clk),
    .D(_01430_),
    .Q(\core.cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16595_ (.CLK(clk),
    .D(_01431_),
    .Q(\core.cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16596_ (.CLK(clk),
    .D(_01432_),
    .Q(\core.cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16597_ (.CLK(clk),
    .D(_01433_),
    .Q(\core.cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16598_ (.CLK(clk),
    .D(_01434_),
    .Q(\core.cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16599_ (.CLK(clk),
    .D(_01435_),
    .Q(\core.cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16600_ (.CLK(clk),
    .D(_01436_),
    .Q(\core.cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16601_ (.CLK(clk),
    .D(_01437_),
    .Q(\core.cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16602_ (.CLK(clk),
    .D(_01438_),
    .Q(\core.cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16603_ (.CLK(clk),
    .D(_01439_),
    .Q(\core.cpuregs[24][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16604_ (.CLK(clk),
    .D(_01440_),
    .Q(\core.cpuregs[24][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16605_ (.CLK(clk),
    .D(_01441_),
    .Q(\core.cpuregs[24][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16606_ (.CLK(clk),
    .D(_01442_),
    .Q(\core.cpuregs[24][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16607_ (.CLK(clk),
    .D(_01443_),
    .Q(\core.cpuregs[24][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16608_ (.CLK(clk),
    .D(_01444_),
    .Q(\core.cpuregs[24][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16609_ (.CLK(clk),
    .D(_01445_),
    .Q(\core.cpuregs[24][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16610_ (.CLK(clk),
    .D(_01446_),
    .Q(\core.cpuregs[24][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16611_ (.CLK(clk),
    .D(_01447_),
    .Q(\core.cpuregs[24][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16612_ (.CLK(clk),
    .D(_01448_),
    .Q(\core.cpuregs[24][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16613_ (.CLK(clk),
    .D(_01449_),
    .Q(\core.cpuregs[24][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16614_ (.CLK(clk),
    .D(_01450_),
    .Q(\core.cpuregs[24][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16615_ (.CLK(clk),
    .D(_01451_),
    .Q(\core.cpuregs[24][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16616_ (.CLK(clk),
    .D(_01452_),
    .Q(\core.cpuregs[24][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16617_ (.CLK(clk),
    .D(_01453_),
    .Q(\core.cpuregs[24][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16618_ (.CLK(clk),
    .D(_01454_),
    .Q(\core.cpuregs[24][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16619_ (.CLK(clk),
    .D(_01455_),
    .Q(\core.cpuregs[24][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16620_ (.CLK(clk),
    .D(_01456_),
    .Q(\core.cpuregs[24][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16621_ (.CLK(clk),
    .D(_01457_),
    .Q(\core.cpuregs[24][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16622_ (.CLK(clk),
    .D(_01458_),
    .Q(\core.cpuregs[24][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16623_ (.CLK(clk),
    .D(_01459_),
    .Q(\core.cpuregs[24][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16624_ (.CLK(clk),
    .D(_01460_),
    .Q(\core.cpuregs[24][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16625_ (.CLK(clk),
    .D(_01461_),
    .Q(\core.cpuregs[24][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16626_ (.CLK(clk),
    .D(_01462_),
    .Q(\core.cpuregs[24][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16627_ (.CLK(clk),
    .D(_01463_),
    .Q(\core.cpuregs[24][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16628_ (.CLK(clk),
    .D(_01464_),
    .Q(\core.cpuregs[24][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16629_ (.CLK(clk),
    .D(_01465_),
    .Q(\core.cpuregs[24][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16630_ (.CLK(clk),
    .D(_01466_),
    .Q(\core.cpuregs[24][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16631_ (.CLK(clk),
    .D(_01467_),
    .Q(\core.cpuregs[24][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16632_ (.CLK(clk),
    .D(_01468_),
    .Q(\core.cpuregs[24][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16633_ (.CLK(clk),
    .D(_01469_),
    .Q(\core.cpuregs[24][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16634_ (.CLK(clk),
    .D(_01470_),
    .Q(\core.cpuregs[24][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16635_ (.CLK(clk),
    .D(_01471_),
    .Q(\core.cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _16636_ (.CLK(clk),
    .D(_01472_),
    .Q(\core.cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _16637_ (.CLK(clk),
    .D(_01473_),
    .Q(\core.cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _16638_ (.CLK(clk),
    .D(_01474_),
    .Q(\core.cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _16639_ (.CLK(clk),
    .D(_01475_),
    .Q(\core.cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _16640_ (.CLK(clk),
    .D(_01476_),
    .Q(\core.cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _16641_ (.CLK(clk),
    .D(_01477_),
    .Q(\core.cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _16642_ (.CLK(clk),
    .D(_01478_),
    .Q(\core.cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _16643_ (.CLK(clk),
    .D(_01479_),
    .Q(\core.cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _16644_ (.CLK(clk),
    .D(_01480_),
    .Q(\core.cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _16645_ (.CLK(clk),
    .D(_01481_),
    .Q(\core.cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _16646_ (.CLK(clk),
    .D(_01482_),
    .Q(\core.cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _16647_ (.CLK(clk),
    .D(_01483_),
    .Q(\core.cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _16648_ (.CLK(clk),
    .D(_01484_),
    .Q(\core.cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _16649_ (.CLK(clk),
    .D(_01485_),
    .Q(\core.cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _16650_ (.CLK(clk),
    .D(_01486_),
    .Q(\core.cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _16651_ (.CLK(clk),
    .D(_01487_),
    .Q(\core.cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _16652_ (.CLK(clk),
    .D(_01488_),
    .Q(\core.cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _16653_ (.CLK(clk),
    .D(_01489_),
    .Q(\core.cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _16654_ (.CLK(clk),
    .D(_01490_),
    .Q(\core.cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _16655_ (.CLK(clk),
    .D(_01491_),
    .Q(\core.cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _16656_ (.CLK(clk),
    .D(_01492_),
    .Q(\core.cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _16657_ (.CLK(clk),
    .D(_01493_),
    .Q(\core.cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _16658_ (.CLK(clk),
    .D(_01494_),
    .Q(\core.cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _16659_ (.CLK(clk),
    .D(_01495_),
    .Q(\core.cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _16660_ (.CLK(clk),
    .D(_01496_),
    .Q(\core.cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _16661_ (.CLK(clk),
    .D(_01497_),
    .Q(\core.cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _16662_ (.CLK(clk),
    .D(_01498_),
    .Q(\core.cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _16663_ (.CLK(clk),
    .D(_01499_),
    .Q(\core.cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _16664_ (.CLK(clk),
    .D(_01500_),
    .Q(\core.cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _16665_ (.CLK(clk),
    .D(_01501_),
    .Q(\core.cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _16666_ (.CLK(clk),
    .D(_01502_),
    .Q(\core.cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _16667_ (.CLK(clk),
    .D(_01503_),
    .Q(\core.instr_lhu ));
 sky130_fd_sc_hd__dfxtp_2 _16668_ (.CLK(clk),
    .D(_01504_),
    .Q(\core.instr_lbu ));
 sky130_fd_sc_hd__dfxtp_2 _16669_ (.CLK(clk),
    .D(_01505_),
    .Q(\core.instr_lw ));
 sky130_fd_sc_hd__dfxtp_2 _16670_ (.CLK(clk),
    .D(_01506_),
    .Q(\core.instr_lh ));
 sky130_fd_sc_hd__dfxtp_2 _16671_ (.CLK(clk),
    .D(_01507_),
    .Q(\core.instr_bgeu ));
 sky130_fd_sc_hd__dfxtp_2 _16672_ (.CLK(clk),
    .D(_01508_),
    .Q(\core.instr_blt ));
 sky130_fd_sc_hd__dfxtp_2 _16673_ (.CLK(clk),
    .D(_00034_),
    .Q(\core.reg_sh[2] ));
 sky130_fd_sc_hd__dfxtp_2 _16674_ (.CLK(clk),
    .D(_00035_),
    .Q(\core.reg_sh[3] ));
 sky130_fd_sc_hd__dfxtp_2 _16675_ (.CLK(clk),
    .D(_00036_),
    .Q(\core.reg_sh[4] ));
 sky130_fd_sc_hd__dfxtp_2 _16676_ (.CLK(clk),
    .D(_01509_),
    .Q(\core.instr_rdinstrh ));
 sky130_fd_sc_hd__dfxtp_2 _16677_ (.CLK(clk),
    .D(_00020_),
    .Q(_00000_));
 sky130_fd_sc_hd__dfxtp_2 _16678_ (.CLK(clk),
    .D(_00021_),
    .Q(_00001_));
 sky130_fd_sc_hd__dfxtp_2 _16679_ (.CLK(clk),
    .D(_00022_),
    .Q(_00002_));
 sky130_fd_sc_hd__dfxtp_2 _16680_ (.CLK(clk),
    .D(_00023_),
    .Q(_00003_));
 sky130_fd_sc_hd__dfxtp_2 _16681_ (.CLK(clk),
    .D(_00024_),
    .Q(_00004_));
 sky130_fd_sc_hd__dfxtp_2 _16682_ (.CLK(clk),
    .D(_01510_),
    .Q(\core.instr_rdinstr ));
 sky130_fd_sc_hd__dfxtp_2 _16683_ (.CLK(clk),
    .D(_01511_),
    .Q(\core.instr_rdcycle ));
 sky130_fd_sc_hd__dfxtp_2 _16684_ (.CLK(clk),
    .D(_01512_),
    .Q(\core.instr_srai ));
 sky130_fd_sc_hd__dfxtp_2 _16685_ (.CLK(clk),
    .D(_01513_),
    .Q(\core.instr_and ));
 sky130_fd_sc_hd__dfxtp_2 _16686_ (.CLK(clk),
    .D(_01514_),
    .Q(\core.instr_or ));
 sky130_fd_sc_hd__dfxtp_2 _16687_ (.CLK(clk),
    .D(_01515_),
    .Q(\core.instr_srl ));
 sky130_fd_sc_hd__dfxtp_2 _16688_ (.CLK(clk),
    .D(_01516_),
    .Q(\core.instr_sltu ));
 sky130_fd_sc_hd__dfxtp_2 _16689_ (.CLK(clk),
    .D(_01517_),
    .Q(\core.instr_slt ));
 sky130_fd_sc_hd__dfxtp_2 _16690_ (.CLK(clk),
    .D(_01518_),
    .Q(\core.instr_sub ));
 sky130_fd_sc_hd__dfxtp_2 _16691_ (.CLK(clk),
    .D(_01519_),
    .Q(\core.instr_slli ));
 sky130_fd_sc_hd__dfxtp_2 _16692_ (.CLK(clk),
    .D(_01520_),
    .Q(\core.instr_sw ));
 sky130_fd_sc_hd__dfxtp_2 _16693_ (.CLK(clk),
    .D(_01521_),
    .Q(\core.instr_andi ));
 sky130_fd_sc_hd__dfxtp_2 _16694_ (.CLK(clk),
    .D(_01522_),
    .Q(\core.instr_xori ));
 sky130_fd_sc_hd__dfxtp_2 _16695_ (.CLK(clk),
    .D(_01523_),
    .Q(\core.instr_addi ));
 sky130_fd_sc_hd__dfxtp_2 _16696_ (.CLK(clk),
    .D(_01524_),
    .Q(\core.instr_sb ));
 sky130_fd_sc_hd__dfxtp_2 _16697_ (.CLK(clk),
    .D(_01525_),
    .Q(\core.mem_do_rdata ));
 sky130_fd_sc_hd__dfxtp_2 _16698_ (.CLK(clk),
    .D(_01526_),
    .Q(\core.mem_do_rinst ));
 sky130_fd_sc_hd__dfxtp_2 _16699_ (.CLK(clk),
    .D(_01527_),
    .Q(\core.mem_do_prefetch ));
 sky130_fd_sc_hd__dfxtp_2 _16700_ (.CLK(clk),
    .D(_01528_),
    .Q(mem_addr[2]));
 sky130_fd_sc_hd__dfxtp_2 _16701_ (.CLK(clk),
    .D(_01529_),
    .Q(mem_addr[3]));
 sky130_fd_sc_hd__dfxtp_2 _16702_ (.CLK(clk),
    .D(_01530_),
    .Q(mem_addr[4]));
 sky130_fd_sc_hd__dfxtp_2 _16703_ (.CLK(clk),
    .D(_01531_),
    .Q(mem_addr[5]));
 sky130_fd_sc_hd__dfxtp_2 _16704_ (.CLK(clk),
    .D(_01532_),
    .Q(mem_addr[6]));
 sky130_fd_sc_hd__dfxtp_2 _16705_ (.CLK(clk),
    .D(_01533_),
    .Q(mem_addr[7]));
 sky130_fd_sc_hd__dfxtp_2 _16706_ (.CLK(clk),
    .D(_01534_),
    .Q(mem_addr[8]));
 sky130_fd_sc_hd__dfxtp_2 _16707_ (.CLK(clk),
    .D(_01535_),
    .Q(mem_addr[9]));
 sky130_fd_sc_hd__dfxtp_2 _16708_ (.CLK(clk),
    .D(_01536_),
    .Q(mem_addr[10]));
 sky130_fd_sc_hd__dfxtp_2 _16709_ (.CLK(clk),
    .D(_01537_),
    .Q(mem_addr[11]));
 sky130_fd_sc_hd__dfxtp_2 _16710_ (.CLK(clk),
    .D(_01538_),
    .Q(mem_addr[12]));
 sky130_fd_sc_hd__dfxtp_2 _16711_ (.CLK(clk),
    .D(_01539_),
    .Q(mem_addr[13]));
 sky130_fd_sc_hd__dfxtp_2 _16712_ (.CLK(clk),
    .D(_01540_),
    .Q(mem_addr[14]));
 sky130_fd_sc_hd__dfxtp_2 _16713_ (.CLK(clk),
    .D(_01541_),
    .Q(mem_addr[15]));
 sky130_fd_sc_hd__dfxtp_2 _16714_ (.CLK(clk),
    .D(_01542_),
    .Q(mem_addr[16]));
 sky130_fd_sc_hd__conb_1 _16715_ (.LO(mem_addr[0]));
 sky130_fd_sc_hd__conb_1 _16716_ (.LO(mem_addr[1]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
endmodule
